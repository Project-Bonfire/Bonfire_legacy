--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated!
-- Here are the parameters:
-- 	 network size x:2
-- 	 network size y:2
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.TB_Package.all;

USE ieee.numeric_std.ALL; 
use IEEE.math_real."ceil";
use IEEE.math_real."log2";

entity tb_network_2x2 is
end tb_network_2x2; 


architecture behavior of tb_network_2x2 is

-- Declaring network component
component network_2x2 is
 generic (DATA_WIDTH: integer := 32; DATA_WIDTH_LV: integer := 11);
port (reset: in  std_logic; 
	clk: in  std_logic; 
	--------------
	RX_L_0: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_0, valid_out_L_0: out std_logic;
	credit_in_L_0, valid_in_L_0: in std_logic;
	TX_L_0: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_1: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_1, valid_out_L_1: out std_logic;
	credit_in_L_1, valid_in_L_1: in std_logic;
	TX_L_1: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_2: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_2, valid_out_L_2: out std_logic;
	credit_in_L_2, valid_in_L_2: in std_logic;
	TX_L_2: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_3: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_3, valid_out_L_3: out std_logic;
	credit_in_L_3, valid_in_L_3: in std_logic;
	TX_L_3: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--fault injector signals
	FI_Add_2_0, FI_Add_0_2: in std_logic_vector(4 downto 0);
	sta0_0_2, sta1_0_2, sta0_2_0, sta1_2_0: in std_logic;

	FI_Add_3_1, FI_Add_1_3: in std_logic_vector(4 downto 0);
	sta0_1_3, sta1_1_3, sta0_3_1, sta1_3_1: in std_logic;

	FI_Add_1_0, FI_Add_0_1: in std_logic_vector(4 downto 0);
	sta0_0_1, sta1_0_1, sta0_1_0, sta1_1_0: in std_logic;

	FI_Add_3_2, FI_Add_2_3: in std_logic_vector(4 downto 0);
	sta0_2_3, sta1_2_3, sta0_3_2, sta1_3_2: in std_logic;

	--------------
    link_faults_0: out std_logic_vector(4 downto 0);
    turn_faults_0: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_0: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_0: in  std_logic_vector(3 downto 0);
    Reconfig_command_0 : in std_logic;

	--------------
    link_faults_1: out std_logic_vector(4 downto 0);
    turn_faults_1: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_1: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_1: in  std_logic_vector(3 downto 0);
    Reconfig_command_1 : in std_logic;

	--------------
    link_faults_2: out std_logic_vector(4 downto 0);
    turn_faults_2: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_2: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_2: in  std_logic_vector(3 downto 0);
    Reconfig_command_2 : in std_logic;

	--------------
    link_faults_3: out std_logic_vector(4 downto 0);
    turn_faults_3: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_3: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_3: in  std_logic_vector(3 downto 0);
    Reconfig_command_3 : in std_logic
            ); 
end component; 
component NoC_Node is
generic( current_address : integer := 0;
         stim_file: string :="code.txt";
         log_file  : string := "output.txt");

port( reset        : in std_logic;
      clk          : in std_logic;

        credit_in : in std_logic;
        valid_out: out std_logic;
        TX: out std_logic_vector(31 downto 0);

        credit_out : out std_logic;
        valid_in: in std_logic;
        RX: in std_logic_vector(31 downto 0);

        link_faults: in std_logic_vector(4 downto 0);
        turn_faults: in std_logic_vector(19 downto 0);

        Rxy_reconf_PE: out  std_logic_vector(7 downto 0);
        Cx_reconf_PE: out  std_logic_vector(3 downto 0);
        Reconfig_command : out std_logic

   );
end component; --component NoC_Node

-- generating bulk signals...
	signal RX_L_0, TX_L_0:  std_logic_vector (31 downto 0);
	signal credit_counter_out_0:  std_logic_vector (1 downto 0);
	signal credit_out_L_0, credit_in_L_0, valid_in_L_0, valid_out_L_0: std_logic;
	signal RX_L_1, TX_L_1:  std_logic_vector (31 downto 0);
	signal credit_counter_out_1:  std_logic_vector (1 downto 0);
	signal credit_out_L_1, credit_in_L_1, valid_in_L_1, valid_out_L_1: std_logic;
	signal RX_L_2, TX_L_2:  std_logic_vector (31 downto 0);
	signal credit_counter_out_2:  std_logic_vector (1 downto 0);
	signal credit_out_L_2, credit_in_L_2, valid_in_L_2, valid_out_L_2: std_logic;
	signal RX_L_3, TX_L_3:  std_logic_vector (31 downto 0);
	signal credit_counter_out_3:  std_logic_vector (1 downto 0);
	signal credit_out_L_3, credit_in_L_3, valid_in_L_3, valid_out_L_3: std_logic;
	--fault injector signals
	signal FI_Add_2_0, FI_Add_0_2: std_logic_vector(integer(ceil(log2(real(31))))-1 downto 0) := (others=>'0');
	signal sta0_0_2, sta1_0_2, sta0_2_0, sta1_2_0: std_logic :='0';

	signal FI_Add_3_1, FI_Add_1_3: std_logic_vector(integer(ceil(log2(real(31))))-1 downto 0) := (others=>'0');
	signal sta0_1_3, sta1_1_3, sta0_3_1, sta1_3_1: std_logic :='0';

	signal FI_Add_1_0, FI_Add_0_1: std_logic_vector(integer(ceil(log2(real(31))))-1 downto 0):= (others=>'0');
	signal sta0_0_1, sta1_0_1, sta0_1_0, sta1_1_0: std_logic :='0';

	signal FI_Add_3_2, FI_Add_2_3: std_logic_vector(integer(ceil(log2(real(31))))-1 downto 0):= (others=>'0');
	signal sta0_2_3, sta1_2_3, sta0_3_2, sta1_3_2: std_logic :='0';

	signal link_faults_0 : std_logic_vector(4 downto 0);
	signal turn_faults_0 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_0 : std_logic_vector(7 downto 0);
	signal Cx_reconf_PE_0 : std_logic_vector(3 downto 0);
	signal Reconfig_command_0 : std_logic;
	signal link_faults_1 : std_logic_vector(4 downto 0);
	signal turn_faults_1 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_1 : std_logic_vector(7 downto 0);
	signal Cx_reconf_PE_1 : std_logic_vector(3 downto 0);
	signal Reconfig_command_1 : std_logic;
	signal link_faults_2 : std_logic_vector(4 downto 0);
	signal turn_faults_2 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_2 : std_logic_vector(7 downto 0);
	signal Cx_reconf_PE_2 : std_logic_vector(3 downto 0);
	signal Reconfig_command_2 : std_logic;
	signal link_faults_3 : std_logic_vector(4 downto 0);
	signal turn_faults_3 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_3 : std_logic_vector(7 downto 0);
	signal Cx_reconf_PE_3 : std_logic_vector(3 downto 0);
	signal Reconfig_command_3 : std_logic;
	--------------

 constant clk_period : time := 1 ns;
signal reset, not_reset, clk: std_logic :='0';

begin

   clk_process :process
   begin
        clk <= '0';
        wait for clk_period/2;   
        clk <= '1';
        wait for clk_period/2; 
   end process;

reset <= '1' after 1 ns;
-- instantiating the network
NoC: network_2x2 generic map (DATA_WIDTH  => 32, DATA_WIDTH_LV => 11)
port map (reset, clk, 
	RX_L_0, credit_out_L_0, valid_out_L_0, credit_in_L_0, valid_in_L_0,  TX_L_0, 
	RX_L_1, credit_out_L_1, valid_out_L_1, credit_in_L_1, valid_in_L_1,  TX_L_1, 
	RX_L_2, credit_out_L_2, valid_out_L_2, credit_in_L_2, valid_in_L_2,  TX_L_2, 
	RX_L_3, credit_out_L_3, valid_out_L_3, credit_in_L_3, valid_in_L_3,  TX_L_3, 
	--fault injector signals
	--FI vertical signals
	FI_Add_2_0, FI_Add_0_2, 
	sta0_0_2, sta1_0_2, sta0_2_0, sta1_2_0, 
	FI_Add_3_1, FI_Add_1_3, 
	sta0_1_3, sta1_1_3, sta0_3_1, sta1_3_1, 
	--FI horizontal signals
	FI_Add_1_0, FI_Add_0_1,
	sta0_0_1, sta1_0_1, sta0_1_0, sta1_1_0, 
	FI_Add_3_2, FI_Add_2_3,
	sta0_2_3, sta1_2_3, sta0_3_2, sta1_3_2, 
	-- should be connected to NI
	link_faults_0, turn_faults_0,	Rxy_reconf_PE_0, Cx_reconf_PE_0, Reconfig_command_0, 
	link_faults_1, turn_faults_1,	Rxy_reconf_PE_1, Cx_reconf_PE_1, Reconfig_command_1, 
	link_faults_2, turn_faults_2,	Rxy_reconf_PE_2, Cx_reconf_PE_2, Reconfig_command_2, 
	link_faults_3, turn_faults_3,	Rxy_reconf_PE_3, Cx_reconf_PE_3, Reconfig_command_3
            ); 
not_reset <= not reset; 

-- connecting the PEs
PE_0: NoC_Node 
generic map( current_address => 0,
	stim_file => "code_0.txt",
	log_file  => "output_0.txt")

port map( not_reset, clk, 

        credit_in => credit_out_L_0, 
        valid_out => valid_in_L_0,
        TX => RX_L_0, 

        credit_out => credit_in_L_0, 
        valid_in => valid_out_L_0,
        RX => TX_L_0,
        link_faults => link_faults_0,
        turn_faults => turn_faults_0,
        Rxy_reconf_PE => Rxy_reconf_PE_0, 
        Cx_reconf_PE => Cx_reconf_PE_0,
        Reconfig_command => Reconfig_command_0
   );
PE_1: NoC_Node 
generic map( current_address => 1,
	stim_file => "code_1.txt",
	log_file  => "output_1.txt")

port map( not_reset, clk, 

        credit_in => credit_out_L_1, 
        valid_out => valid_in_L_1,
        TX => RX_L_1, 

        credit_out => credit_in_L_1, 
        valid_in => valid_out_L_1,
        RX => TX_L_1,
        link_faults => link_faults_1,
        turn_faults => turn_faults_1,
        Rxy_reconf_PE => Rxy_reconf_PE_1, 
        Cx_reconf_PE => Cx_reconf_PE_1,
        Reconfig_command => Reconfig_command_1
   );
PE_2: NoC_Node 
generic map( current_address => 2,
	stim_file => "code_2.txt",
	log_file  => "output_2.txt")

port map( not_reset, clk, 

        credit_in => credit_out_L_2, 
        valid_out => valid_in_L_2,
        TX => RX_L_2, 

        credit_out => credit_in_L_2, 
        valid_in => valid_out_L_2,
        RX => TX_L_2,
        link_faults => link_faults_2,
        turn_faults => turn_faults_2,
        Rxy_reconf_PE => Rxy_reconf_PE_2, 
        Cx_reconf_PE => Cx_reconf_PE_2,
        Reconfig_command => Reconfig_command_2
   );
PE_3: NoC_Node 
generic map( current_address => 3,
	stim_file => "code_3.txt",
	log_file  => "output_3.txt")

port map( not_reset, clk, 

        credit_in => credit_out_L_3, 
        valid_out => valid_in_L_3,
        TX => RX_L_3, 

        credit_out => credit_in_L_3, 
        valid_in => valid_out_L_3,
        RX => TX_L_3,
        link_faults => link_faults_3,
        turn_faults => turn_faults_3,
        Rxy_reconf_PE => Rxy_reconf_PE_3, 
        Cx_reconf_PE => Cx_reconf_PE_3,
        Reconfig_command => Reconfig_command_3
   );

-- connecting the fault generators
gen_fault(sta0_1_0, sta1_1_0, FI_Add_1_0, 56,1138666221,1960809222);
gen_fault(sta0_0_1, sta1_0_1, FI_Add_0_1, 64,751500117,1520623220);
gen_fault(sta0_2_0, sta1_2_0, FI_Add_2_0, 70,1730004934,1255590821);
gen_fault(sta0_0_2, sta1_0_2, FI_Add_0_2, 45,332821241,1061603537);
gen_fault(sta0_3_1, sta1_3_1, FI_Add_3_1, 53,750959745,841254867);
gen_fault(sta0_1_3, sta1_1_3, FI_Add_1_3, 46,1831451386,1574401837);
gen_fault(sta0_3_2, sta1_3_2, FI_Add_3_2, 57,929911280,1401056219);
gen_fault(sta0_2_3, sta1_2_3, FI_Add_2_3, 59,322054547,1380824540);


end;
