--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated!
-- Here are the parameters:
-- 	 network size x: 2
-- 	 network size y: 2
-- 	 Data width: 32
-- 	 Parity: False
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.numeric_std.ALL;
use work.component_pack.all;

entity network_2x2_with_PE is
 generic (DATA_WIDTH: integer := 32;
          DATA_WIDTH_LV: integer := 11;
          memory_type : string :=
            "TRI_PORT_X"
           --   "DUAL_PORT_"
           --   "ALTERA_LPM"
           --   "XILINX_16X"
      );

port (reset: in  std_logic;
      clk: in  std_logic;

      -- IJTAG network for fault injection and checker status monitoring
      TCK         : in std_logic;
      RST         : in std_logic;
      SEL         : in std_logic;
      SI          : in std_logic;
      SE          : in std_logic;
      UE          : in std_logic;
      CE          : in std_logic;
      SO          : out std_logic;
      toF         : out std_logic;
      toC         : out std_logic;

      -- GPIO for Node 0
      GPIO_out: out  std_logic_vector(15 downto 0);
      GPIO_in: in  std_logic_vector(21 downto 0);

      -- UART for all Plasmas
      uart_write_0  : out std_logic;
      uart_read_0   : in std_logic;
      uart_write_1  : out std_logic;
      uart_read_1   : in std_logic;
      uart_write_2  : out std_logic;
      uart_read_2   : in std_logic;
      uart_write_3  : out std_logic;
      uart_read_3   : in std_logic;

      -- Monitor connections
      temperature_control   : out std_logic_vector(3 downto 0);
      temperature_data      : in std_logic_vector(12 downto 0);
      iddt_control          : out std_logic_vector(2 downto 0);
      iddt_data             : in std_logic_vector(12 downto 0);
      slack_control         : out std_logic_vector(2 downto 0);
      slack_data            : in std_logic_vector(31 downto 0);
      voltage_control       : out std_logic_vector(2 downto 0);
      voltage_data          : in std_logic_vector(31 downto 0)
    );

end network_2x2_with_PE;


architecture behavior of network_2x2_with_PE is

constant path : string(1 to 12) := "Testbenches/"; --uncomment this if you are SIMULATING in MODELSIM, or if you're synthesizing.
-- constant path : string(positive range <>) := "/home/tsotne/ownCloud/git/Bonfire_sim/Bonfire/RTL/Chip_Designs/IMMORTAL_Chip_2017/Testbenches/"; --used only for Vivado similation. Tsotnes PC.

    component immortal_sensor_IJTAG_interface is
    Port ( -- Scan Interface  client --------------
            TCK         : in std_logic;
            RST         : in std_logic;
            SEL         : in std_logic;
            SI          : in std_logic;
            SE          : in std_logic;
            UE          : in std_logic;
            CE          : in std_logic;
            SO          : out std_logic;
            toF         : out std_logic;
            toC         : out std_logic;

            -- Monitor connections
            temperature_control   : out std_logic_vector(3 downto 0);
            temperature_data      : in std_logic_vector(12 downto 0);
            iddt_control          : out std_logic_vector(2 downto 0);
            iddt_data             : in std_logic_vector(12 downto 0);
            slack_control         : out std_logic_vector(2 downto 0);
            slack_data            : in std_logic_vector(31 downto 0);
            voltage_control       : out std_logic_vector(2 downto 0);
            voltage_data          : in std_logic_vector(31 downto 0));
    end component;

-- Declaring network component

-- Declaring NoC_Node component (with Plasma, RAM, NI and UART)


-- generating bulk signals...
    signal RX_L_0, TX_L_0:  std_logic_vector (31 downto 0);
    signal credit_counter_out_0:  std_logic_vector (1 downto 0);
    signal credit_out_L_0, credit_in_L_0, valid_in_L_0, valid_out_L_0: std_logic;
    signal RX_L_1, TX_L_1:  std_logic_vector (31 downto 0);
    signal credit_counter_out_1:  std_logic_vector (1 downto 0);
    signal credit_out_L_1, credit_in_L_1, valid_in_L_1, valid_out_L_1: std_logic;
    signal RX_L_2, TX_L_2:  std_logic_vector (31 downto 0);
    signal credit_counter_out_2:  std_logic_vector (1 downto 0);
    signal credit_out_L_2, credit_in_L_2, valid_in_L_2, valid_out_L_2: std_logic;
    signal RX_L_3, TX_L_3:  std_logic_vector (31 downto 0);
    signal credit_counter_out_3:  std_logic_vector (1 downto 0);
    signal credit_out_L_3, credit_in_L_3, valid_in_L_3, valid_out_L_3: std_logic;

    -- NI testing signals
    --------------
    --signal Rxy_reconf: std_logic_vector (7 downto 0) := "01111101";
    --signal Reconfig: std_logic := '0';
    --------------

    signal not_reset: std_logic;

    signal link_faults_0, link_faults_1, link_faults_2, link_faults_3   : std_logic_vector(4 downto 0);
    signal turn_faults_0, turn_faults_1, turn_faults_2, turn_faults_3   : std_logic_vector(19 downto 0);
    signal Rxy_reconf_PE_0, Rxy_reconf_PE_1,Rxy_reconf_PE_2, Rxy_reconf_PE_3   : std_logic_vector(7 downto 0);
    signal Cx_reconf_PE_0, Cx_reconf_PE_1, Cx_reconf_PE_2, Cx_reconf_PE_3 : std_logic_vector(3 downto 0);
    signal Reconfig_command_0, Reconfig_command_1, Reconfig_command_2, Reconfig_command_3 : std_logic;

    signal GPIO_out_FF_in, GPIO_out_FF : std_logic_vector(15 downto 0);
    signal UART_0_W_in, UART_0_W_out, UART_0_R_in, UART_0_R_out : std_logic;
    signal UART_1_W_in, UART_1_W_out, UART_1_R_in, UART_1_R_out : std_logic;
    signal UART_2_W_in, UART_2_W_out, UART_2_R_in, UART_2_R_out : std_logic;
    signal UART_3_W_in, UART_3_W_out, UART_3_R_in, UART_3_R_out : std_logic;

    signal SO_NoC , SO_sensors  : std_logic;
    signal toF_NoC, toF_sensors : std_logic;
    signal toC_NoC, toC_sensors : std_logic;

begin

-- instantiating the network
NoC: network_2x2 generic map (DATA_WIDTH  => 32, DATA_WIDTH_LV => 11)
port map (reset, clk,
    RX_L_0, credit_out_L_0, valid_out_L_0, credit_in_L_0, valid_in_L_0,  TX_L_0,
    RX_L_1, credit_out_L_1, valid_out_L_1, credit_in_L_1, valid_in_L_1,  TX_L_1,
    RX_L_2, credit_out_L_2, valid_out_L_2, credit_in_L_2, valid_in_L_2,  TX_L_2,
    RX_L_3, credit_out_L_3, valid_out_L_3, credit_in_L_3, valid_in_L_3,  TX_L_3,
    link_faults_0, turn_faults_0, Rxy_reconf_PE_0, Cx_reconf_PE_0, Reconfig_command_0,
    link_faults_1, turn_faults_1, Rxy_reconf_PE_1, Cx_reconf_PE_1, Reconfig_command_1,
    link_faults_2, turn_faults_2, Rxy_reconf_PE_2, Cx_reconf_PE_2, Reconfig_command_2,
    link_faults_3, turn_faults_3, Rxy_reconf_PE_3, Cx_reconf_PE_3, Reconfig_command_3,
    TCK, RST, SEL, SI, SE, UE, CE, SO_NoC, toF_NoC, toC_NoC
    );

toF <= toF_NoC or toF_sensors;
toC <= toC_NoC and toC_sensors;
SO <= SO_sensors;

immortal_sensor_IJTAG_interface: immortal_sensor_IJTAG_interface
    port map (
    TCK => TCK,
    RST => RST,
    SEL => SEL,
    SI  => SO_NoC,
    SE  => SE,
    UE  => UE,
    CE  => CE,
    SO  => SO_sensors,
    toF => toF_sensors,
    toC => toC_sensors,

    temperature_control => temperature_control,
    temperature_data    => temperature_data,
    iddt_control        => iddt_control,
    iddt_data           => iddt_data,
    slack_control       => slack_control,
    slack_data          => slack_data,
    voltage_control     => voltage_control,
    voltage_data        => voltage_data
  );


process (not_reset, clk)
begin
  if not_reset = '1' then
      GPIO_out_FF <= (others => '0');

      UART_0_W_out <= '0';
      UART_1_W_out <= '0';
      UART_2_W_out <= '0';
      UART_3_W_out <= '0';

      UART_0_R_out <= '0';
      UART_1_R_out <= '0';
      UART_2_R_out <= '0';
      UART_3_R_out <= '0';

  elsif clk'event and clk = '1' then
      GPIO_out_FF <= GPIO_out_FF_in;

      UART_0_W_out <= UART_0_W_in;
      UART_1_W_out <= UART_1_W_in;
      UART_2_W_out <= UART_2_W_in;
      UART_3_W_out <= UART_3_W_in;

      UART_0_R_out <= UART_0_R_in;
      UART_1_R_out <= UART_1_R_in;
      UART_2_R_out <= UART_2_R_in;
      UART_3_R_out <= UART_3_R_in;
  end if;
end process;


GPIO_out <=  GPIO_out_FF;

uart_write_0 <= UART_0_W_out;
uart_write_1 <= UART_1_W_out;
uart_write_2 <= UART_2_W_out;
uart_write_3 <= UART_3_W_out;

UART_0_R_in <= uart_read_0;
UART_1_R_in <= uart_read_1;
UART_2_R_in <= uart_read_2;
UART_3_R_in <= uart_read_3;

not_reset <= not reset;

-- instantiating and connecting the PEs
PE_0: NoC_Node
generic map( current_address => 0,
    stim_file => path & "code_0.txt",
    log_file  => path & "output_0.txt",
    memory_type => memory_type)

port map( not_reset, clk,
        uart_read         => UART_0_R_out,
        uart_write        => UART_0_W_in,
        credit_in => credit_out_L_0,
        valid_out => valid_in_L_0,
        TX => RX_L_0,

        credit_out => credit_in_L_0,
        valid_in => valid_out_L_0,
        RX => TX_L_0,
        link_faults         => link_faults_0,
        turn_faults         => turn_faults_0,
        Rxy_reconf_PE       => Rxy_reconf_PE_0,
        Cx_reconf_PE        => Cx_reconf_PE_0,
        Reconfig_command    => Reconfig_command_0,

        GPIO_out            => GPIO_out_FF_in,
        GPIO_in             => GPIO_in
   );

PE_1: NoC_Node
generic map( current_address => 1,
    stim_file => path & "code_1.txt",
    log_file  => path & "output_1.txt",
    memory_type => memory_type)

port map( not_reset, clk,
        uart_read         => UART_1_R_out,
        uart_write        => UART_1_W_in,

        credit_in => credit_out_L_1,
        valid_out => valid_in_L_1,
        TX => RX_L_1,

        credit_out => credit_in_L_1,
        valid_in => valid_out_L_1,
        RX => TX_L_1,
        link_faults         => link_faults_1,
        turn_faults         => turn_faults_1,
        Rxy_reconf_PE       => Rxy_reconf_PE_1,
        Cx_reconf_PE        => Cx_reconf_PE_1,
        Reconfig_command    => Reconfig_command_1,

        GPIO_out            => open,
        GPIO_in             => (others => '0')
   );

PE_2: NoC_Node
generic map( current_address => 2,
    stim_file => path & "code_2.txt",
    log_file  => path & "output_2.txt",
    memory_type => memory_type)

port map( not_reset, clk,
        uart_read         => UART_2_R_out,
        uart_write        => UART_2_W_in,

        credit_in => credit_out_L_2,
        valid_out => valid_in_L_2,
        TX => RX_L_2,

        credit_out => credit_in_L_2,
        valid_in => valid_out_L_2,
        RX => TX_L_2,
        link_faults         => link_faults_2,
        turn_faults         => turn_faults_2,
        Rxy_reconf_PE       => Rxy_reconf_PE_2,
        Cx_reconf_PE        => Cx_reconf_PE_2,
        Reconfig_command    => Reconfig_command_2,

        GPIO_out            => open,
        GPIO_in             => (others => '0')
   );

PE_3: NoC_Node
generic map( current_address => 3,
    stim_file => path & "code_3.txt",
    log_file  => path & "output_3.txt",
    memory_type => memory_type)

port map( not_reset, clk,
        uart_read         => UART_3_R_out,
        uart_write        => UART_3_W_in,

        credit_in => credit_out_L_3,
        valid_out => valid_in_L_3,
        TX => RX_L_3,

        credit_out => credit_in_L_3,
        valid_in => valid_out_L_3,
        RX => TX_L_3,
        link_faults         => link_faults_3,
        turn_faults         => turn_faults_3,
        Rxy_reconf_PE       => Rxy_reconf_PE_3,
        Cx_reconf_PE        => Cx_reconf_PE_3,
        Reconfig_command    => Reconfig_command_3,

        GPIO_out            => open,
        GPIO_in             => (others => '0')
   );



end;
