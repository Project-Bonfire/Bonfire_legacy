--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated Please do not change!
-- Here are the parameters:
-- 	 network size x:2
-- 	 network size y:2
-- 	 data width:32-- 	 traffic pattern:------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--use work.TB_Package.all;

USE ieee.numeric_std.ALL;
--use IEEE.math_real."ceil";
--use IEEE.math_real."log2";

entity tb_network_2x2 is
end tb_network_2x2;


architecture behavior of tb_network_2x2 is

-- Declaring network component
component network_2x2_with_PE is
 generic (DATA_WIDTH: integer := 32; DATA_WIDTH_LV: integer := 11);
port (reset: in  std_logic;
      clk: in  std_logic;

      -- IJTAG network for fault injection and checker status monitoring
      TCK         : in std_logic;
      RST         : in std_logic;
      SEL         : in std_logic;
      SI          : in std_logic;
      SE          : in std_logic;
      UE          : in std_logic;
      CE          : in std_logic;
      SO          : out std_logic;
      toF         : out std_logic;
      toC         : out std_logic; 
 
      -- GPIO for Node 0
      GPIO_out: out  std_logic_vector(15 downto 0);
      GPIO_in: in  std_logic_vector(21 downto 0);
           -- UART for all Plasmas
      uart_write_0  : out std_logic;
      uart_read_0   : in std_logic;
      uart_write_1  : out std_logic;
      uart_read_1   : in std_logic;
      uart_write_2  : out std_logic;
      uart_read_2   : in std_logic;
      uart_write_3  : out std_logic;
      uart_read_3   : in std_logic
    );
end component; 

	  constant clk_period : time := 10 ns;
	  constant tck_period : time := 100 ns;
    constant HALF_SEPARATOR : time := 2*tck_period;
    constant FULL_SEPARATOR : time := 8*tck_period;

	  signal reset, not_reset, clk: std_logic :='0';

    signal TCK, RST, SEL, SI, SE, UE, CE, SO, toF, toC : std_logic := '0';

    -- GPIO
    signal PE_0_GPIO_out : std_logic_vector(15 downto 0);
    signal PE_0_GPIO_in : std_logic_vector(21 downto 0) := (others => '1');
    signal uart_write_0,  uart_write_1, uart_write_2, uart_write_3: std_logic;
    signal uart_read_0,   uart_read_1,  uart_read_2,  uart_read_3: std_logic;
begin

  clk_process :process
  begin
      clk <= '0';
      wait for clk_period/2;
      clk <= '1';
      wait for clk_period/2;
  end process;

  ijtag_shift_proc: process

       -- Generate a number of TCK ticks
    procedure tck_tick (number_of_tick : in positive) is
    begin
      for i in 1 to number_of_tick loop
        TCK <= '0';
        wait for TCK_period/2;
        TCK <= '1';
        wait for TCK_period/2;
      end loop;
    end procedure tck_tick;
    
    procedure tck_halftick_high is
    begin
      TCK <= '1';
      wait for TCK_period/2;
    end procedure tck_halftick_high;
             
    procedure tck_halftick_low is
    begin
      TCK <= '0';
      wait for TCK_period/2;
    end procedure tck_halftick_low;

     -- Shifts in specified data (Capture -> Shift -> Update)
    procedure shift_data (data : in std_logic_vector) is
    begin
       -- Capture phase
      --CE <= '1';
      --tck_tick(1);
      --CE <= '0';
        -- Shift phase
      SE <= '1';
      for i in data'range loop
         SI <= data(i);
         tck_tick(1);
      end loop;
      SE <= '0';
      -- Update phase
      UE <= '1';
      tck_tick(1);
      tck_halftick_low;
      UE <= '0';
      tck_halftick_high;
    end procedure shift_data;

          -- Returns all zeroes std_logic_vector of specified size
    function all_zeroes (number_of_zeroes : in positive) return std_logic_vector is
      variable zero_array : std_logic_vector(0 to number_of_zeroes-1);
    begin
      for i in zero_array'range loop
       zero_array(i) := '0';
      end loop;
      return zero_array;
    end function all_zeroes;

  begin

            -- Reset iJTAG chain and Instruments
    RST <= '1';
    wait for tck_period;
    RST <= '0';
    SEL <= '1';
    tck_tick(4);

    --shift_data("0001000000000000"); -- open sib3
    shift_data("0001"&"0000"&"0000"&"0000"); -- open sib3

    tck_tick(4);

    -- 130 bits in total (for chains)
    -- Inject fault in the bit with location 0 of L, N, and W FIFOs , L, N, and W LBDRs , L, N, E, W and S Arbiter_ins and Arbiter_outs and Allocator logic  in Router 3 (SE)
    --shift_data("0000"  & "000000001"     &      "0000001"&"0000001"&"0000001"&"0000001"&"0000001"      &     "0000001"&"0000001"&"0000001"&"0000001"&"0000001"       &"000000001"&"000000001"&"000000001"      &    "00000001"&"00000001"&"00000001"&all_zeroes(12)); --close sib3, shift 1 into the last bit of fault injection register, close other sibs.

    -- Inject fault in the bit with location 0 of L FIFO in Router 3 (SE)
    shift_data("0001"&"0000"&"0001"&"0000"&"0000"&"0000"); --keep sib3 opened, open sib3inj
    shift_data("0001"&"0001"&"0000"& "000000001"     &      "0000001"&"0000001"&"0000001"&"0000001"&"0000001"      &     "0000001"&"0000001"&"0000001"&"0000001"&"0000001"       &"000000001"&"000000001"&"000000001"      &    "00000001"&"00000001"&"00000001"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    shift_data("0001"&"0000"&"1111111111111111111111111"&"0001"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    shift_data("0000"&"0000"&"0000"& "000000001"     &      "0000001"&"0000001"&"0000001"&"0000001"&"0000001"      &     "0000001"&"0000001"&"0000001"&"0000001"&"0000001"       &"000000001"&"000000001"&"000000001"      &    "00000001"&"00000001"&"00000001"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    tck_tick(4);

    shift_data("0001"&"0000"&"0000"&"0000"); -- open sib3

    -- Inject fault in the bit with location 1 of L FIFO in Router 3 (SE)
    shift_data("0001"&"0000"&"0001"&"0000"&"0000"&"0000"); --keep sib3 opened, open sib3inj
    shift_data("0001"&"0001"&"0000"& "000000101"     &      "0000101"&"0000101"&"0000101"&"0000101"&"0000101"      &     "0000101"&"0000101"&"0000101"&"0000101"&"0000101"       &"000000101"&"000000101"&"000000101"      &    "00000101"&"00000101"&"00000101"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    shift_data("0001"&"0000"&"1111111111111111111111111"&"0001"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    shift_data("0000"&"0000"&"0000"& "000000001"     &      "0000101"&"0000101"&"0000101"&"0000101"&"0000101"      &     "0000101"&"0000101"&"0000101"&"0000101"&"0000101"       &"000000101"&"000000101"&"000000101"      &    "00000101"&"00000101"&"00000101"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    tck_tick(4);

    shift_data("0001"&"0000"&"0000"&"0000"); -- open sib3

    -- Inject fault in the bit with location 2 of L FIFO in Router 3 (SE)
    shift_data("0001"&"0000"&"0001"&"0000"&"0000"&"0000"); --keep sib3 opened, open sib3inj
    shift_data("0001"&"0001"&"0000"& "000000001"     &      "0001001"&"0001001"&"0001001"&"0001001"&"0001001"      &     "0001001"&"0001001"&"0001001"&"0001001"&"0001001"       &"000001001"&"000001001"&"000001001"      &    "00001001"&"00001001"&"00001001"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    shift_data("0001"&"0000"&"1111111111111111111111111"&"0001"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    shift_data("0000"&"0000"&"0000"& "000000001"     &      "0001001"&"0001001"&"0001001"&"0001001"&"0001001"      &     "0001001"&"0001001"&"0001001"&"0001001"&"0001001"       &"000001001"&"000001001"&"000001001"      &    "00001001"&"00001001"&"00001001"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    tck_tick(4);

    shift_data("0001"&"0000"&"0000"&"0000"); -- open sib3

    -- Inject fault in the bit with location 3 of L FIFO in Router 3 (SE)
    shift_data("0001"&"0000"&"0001"&"0000"&"0000"&"0000"); --keep sib3 opened, open sib3inj
    shift_data("0001"&"0001"&"0000"& "000000001"     &      "0001101"&"0001101"&"0001101"&"0001101"&"0001101"      &     "0001101"&"0001101"&"0001101"&"0001101"&"0001101"       &"000001101"&"000001101"&"000001101"      &    "00001101"&"00001101"&"00001101"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    shift_data("0001"&"0000"&"1111111111111111111111111"&"0001"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    shift_data("0000"&"0000"&"0000"& "000000001"     &      "0001101"&"0001101"&"0001101"&"0001101"&"0001101"      &     "0001101"&"0001101"&"0001101"&"0001101"&"0001101"       &"000001101"&"000001101"&"000001101"      &    "00001101"&"00001101"&"00001101"&all_zeroes(12)); --close sib3, leave sib3sta closed, shift into fault injection register, close other sibs.
    tck_tick(4);

    wait;

end process;

-- Added for IJTAG

reset <= '1' after 3 ns;

-- instantiating the top module for the network
NoC_top: network_2x2_with_PE generic map (DATA_WIDTH  => 32, DATA_WIDTH_LV => 11)
port map (reset, clk,
	        TCK, RST, SEL, SI, SE, UE, CE, SO, toF, toC, 
          PE_0_GPIO_out, PE_0_GPIO_in, 
          uart_write_0, uart_read_0, 
          uart_write_1, uart_read_1, 
          uart_write_2, uart_read_2, 
          uart_write_3, uart_read_3
         );

end;
