--Copyright (C) 2016 Siavoosh Payandeh Azad

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Arbiter is
    port (  reset: in  std_logic;
            clk: in  std_logic;
            Req_N, Req_E, Req_W, Req_S, Req_L:in std_logic; -- From LBDR modules
            DCTS: in std_logic; -- Getting the CTS signal from the input FIFO of the next router/NI (for hand-shaking)
            Grant_N, Grant_E, Grant_W, Grant_S, Grant_L:out std_logic; -- Grants given to LBDR requests (encoded as one-hot)
            Xbar_sel : out std_logic_vector(4 downto 0); -- select lines for XBAR
            RTS: out std_logic -- Valid output which is sent to the next router/NI to specify that the data on the output port is valid
            );
end;

architecture behavior of Arbiter is
--                                                                        next
--                                     Arbiter                        router or NI
--                     --- ---------------------------- ----          ----
--   from LBDR  --->  |Req(s)                           RTS | -----> |DRTS
--    To FIFO   <---  |Grant(s)                         DCTS| <----- |CTS
--    to XBAR   <---  |Xbar_sel                             |        | 
--                     --- ---------------------------- ----          ----

TYPE STATE_TYPE IS (IDLE, North, East, West, South, Local);
SIGNAL state,next_state   : STATE_TYPE := IDLE;

SIGNAL RTS_FF: std_logic;

begin
		-- process for updating the state of arbiter's FSM, also setting RTS based on the state (if Grant is given or not)
        process(clk,reset)begin
            if reset = '0' then
                state<=IDLE;
                RTS_FF <= '0';
            elsif clk'event and clk = '1' then
                -- no grant given yet, it might be that there is no request to 
                -- arbiter or request is there, but the next router's/NI's FIFO is full
                if next_state = IDLE then 
                    RTS_FF <= '0';
                -- if there was a grant given to one of the inputs, 
                -- tell the next router/NI that the output data is valid
                else 
                    if RTS_ff = '1' and DCTS = '1' then
                        RTS_FF <= '0';
                    else 
                        RTS_FF <= '1';
                    end if;
                end if ;
                state <= next_state;
             end if;
	end process;

    RTS <= RTS_FF;

        -- sets the grants using round robin 
        -- the order is   L --> N --> E --> W --> S 
        process(state, Req_N, Req_E, Req_W, Req_S, Req_L, DCTS)begin
            Grant_N <= '0';
            Grant_E <= '0';
            Grant_W <= '0';
            Grant_S <= '0';
            Grant_L <= '0';
            case(state) is
                when IDLE =>
                    Xbar_sel<= "00000"; 
                    
                    If Req_L = '1' then
                        next_state <= Local;
                    elsif Req_N = '1' then
                        next_state <= North;         
                    elsif Req_E = '1' then
                        next_state <= East;
                    elsif Req_W = '1' then
                        next_state <= West;
                    elsif Req_S = '1' then
                        next_state <= South;
                    else
                        next_state <= IDLE;
                    end if;    
                    
                when North =>
                    Grant_N <= DCTS;

                    Xbar_sel<= "00001";
                    
                    If Req_N = '1' then 
                        next_state <= North; 
                    elsif Req_E = '1' then
                        next_state <= East;
                    elsif Req_W = '1' then
                        next_state <= West;
                    elsif Req_S = '1' then
                        next_state <= South;
                    elsif Req_L = '1' then
                        next_state <= Local;
                    else
                        next_state <= IDLE; 
                    end if;
                    
                when East =>
                    Grant_E <= DCTS;
                    Xbar_sel<= "00010";
                    
                    If Req_E = '1' then 
                        next_state <= East; 
                    elsif Req_W = '1' then
                        next_state <= West;
                    elsif Req_S = '1' then
                        next_state <= South;
                    elsif Req_L = '1' then
                        next_state <= Local;
                    elsif Req_N = '1' then
                        next_state <= North;
                    else
                        next_state <= IDLE; 
                    end if;
                    
                when West =>
                    Grant_W <= DCTS;
                    Xbar_sel<= "00100";
                    
                    If Req_W = '1' then
                        next_state <= West; 
                    elsif Req_S = '1' then
                        next_state <= South;
                    elsif Req_L = '1' then
                        next_state <= Local;
                    elsif Req_N = '1' then
                        next_state <= North;
                    elsif Req_E = '1' then
                        next_state <= East;
                    else
                        next_state <= IDLE; 
                    end if;
                    
                when South =>
                    Grant_S <= DCTS;
                    Xbar_sel<= "01000";
                    
                    If Req_S = '1' then 
                        next_state <= South; 
                    elsif Req_L = '1' then
                        next_state <= Local;
                    elsif Req_N = '1' then
                        next_state <= North;
                    elsif Req_E = '1' then
                        next_state <= East;
                    elsif Req_W = '1' then
                        next_state <= West;
                    else
                        next_state <= IDLE; 
                    end if;
                    
                when Local =>
                    Grant_L <= DCTS;
                    Xbar_sel<= "10000";
                    
                    If Req_L = '1' then
                        next_state <= Local; 
                    elsif Req_N = '1' then
                        next_state <= North;         
                    elsif Req_E = '1' then
                        next_state <= East;
                    elsif Req_W = '1' then
                        next_state <= West;
                    elsif Req_S = '1' then
                        next_state <= South;
                    else
                        next_state <= IDLE; 
                    end if;
                when others =>  
                    null;
            end case ;
        end process;

end;