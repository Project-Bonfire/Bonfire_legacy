--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated Please do not change!
-- Here are the parameters:
-- 	 network size x:2
-- 	 network size y:2
-- 	 data width:32-- 	 traffic pattern:------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--use work.TB_Package.all;

USE ieee.numeric_std.ALL;
--use IEEE.math_real."ceil";
--use IEEE.math_real."log2";

entity mem_wrap_tb is
end mem_wrap_tb;


architecture behavior of mem_wrap_tb is

-- Declaring network component
 

	  constant clk_period : time := 10 ns;

  signal clk, reset, enable: std_logic := '0';
  signal write_byte_enable: std_logic_vector(3 downto 0);
  signal address: std_logic_vector(31 downto 2);
  signal data_write, data_read:  std_logic_vector(31 downto 0);

  component ram is
  generic(memory_type : string := "DEFAULT";
           stim_file: string :="code.txt");
  port(clk               : in std_logic;
        reset             : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
  end component; --entity ram

begin

  clk_process :process
  begin
      clk <= '0';
      wait for clk_period/2;
      clk <= '1';
      wait for clk_period/2;
  end process;

reset <= '1' after clk_period;

 ram_unit: ram port map(clk, reset, enable, write_byte_enable, address, data_write, data_read);

 process(clk)
 variable counter: integer := 0;
 begin
  if reset = '0' then 
    counter := 0;
    enable <= '0'; 
    write_byte_enable <= "0000";
    address <=  (others => '0');
    data_write <= (others => '0');
  elsif falling_edge(clk) then 
    if counter < 10 then
      enable <= '1'; 
      address <=  address + 1;
      write_byte_enable <= "1111";
      data_write <= data_write + 1;
      counter := counter +1;
    else
      if counter < 20 then
        address <=  address - 1;
        enable <= '1'; 
        write_byte_enable <= "0000";
        counter := counter +1;
      else
        enable <= '0';
      end if;
    end if;
  end if;
 end process;
end;
