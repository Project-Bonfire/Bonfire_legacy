--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated!
-- Here are the parameters:
-- 	 network size x:4
-- 	 network size y:4
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.TB_package.all;

entity tb_network_4x4 is
end tb_network_4x4; 


architecture behavior of tb_network_4x4 is

-- Declaring network component
component network_4x4 is
 generic (DATA_WIDTH: integer := 32);
port (reset: in  std_logic; 
	clk: in  std_logic; 
	--------------
	RX_L_0: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_0, CTS_L_0: out std_logic;
	DRTS_L_0, DCTS_L_0: in std_logic;
	TX_L_0: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_1: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_1, CTS_L_1: out std_logic;
	DRTS_L_1, DCTS_L_1: in std_logic;
	TX_L_1: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_2: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_2, CTS_L_2: out std_logic;
	DRTS_L_2, DCTS_L_2: in std_logic;
	TX_L_2: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_3: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_3, CTS_L_3: out std_logic;
	DRTS_L_3, DCTS_L_3: in std_logic;
	TX_L_3: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_4: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_4, CTS_L_4: out std_logic;
	DRTS_L_4, DCTS_L_4: in std_logic;
	TX_L_4: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_5: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_5, CTS_L_5: out std_logic;
	DRTS_L_5, DCTS_L_5: in std_logic;
	TX_L_5: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_6: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_6, CTS_L_6: out std_logic;
	DRTS_L_6, DCTS_L_6: in std_logic;
	TX_L_6: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_7: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_7, CTS_L_7: out std_logic;
	DRTS_L_7, DCTS_L_7: in std_logic;
	TX_L_7: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_8: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_8, CTS_L_8: out std_logic;
	DRTS_L_8, DCTS_L_8: in std_logic;
	TX_L_8: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_9: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_9, CTS_L_9: out std_logic;
	DRTS_L_9, DCTS_L_9: in std_logic;
	TX_L_9: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_10: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_10, CTS_L_10: out std_logic;
	DRTS_L_10, DCTS_L_10: in std_logic;
	TX_L_10: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_11: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_11, CTS_L_11: out std_logic;
	DRTS_L_11, DCTS_L_11: in std_logic;
	TX_L_11: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_12: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_12, CTS_L_12: out std_logic;
	DRTS_L_12, DCTS_L_12: in std_logic;
	TX_L_12: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_13: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_13, CTS_L_13: out std_logic;
	DRTS_L_13, DCTS_L_13: in std_logic;
	TX_L_13: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_14: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_14, CTS_L_14: out std_logic;
	DRTS_L_14, DCTS_L_14: in std_logic;
	TX_L_14: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_15: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_15, CTS_L_15: out std_logic;
	DRTS_L_15, DCTS_L_15: in std_logic;
	TX_L_15: out std_logic_vector (DATA_WIDTH-1 downto 0)
            ); 
end component; 

-- generating bulk signals...
	signal RX_L_0, TX_L_0:  std_logic_vector (31 downto 0);
	signal RTS_L_0, DRTS_L_0, CTS_L_0, DCTS_L_0: std_logic;
	--------------
	signal RX_L_1, TX_L_1:  std_logic_vector (31 downto 0);
	signal RTS_L_1, DRTS_L_1, CTS_L_1, DCTS_L_1: std_logic;
	--------------
	signal RX_L_2, TX_L_2:  std_logic_vector (31 downto 0);
	signal RTS_L_2, DRTS_L_2, CTS_L_2, DCTS_L_2: std_logic;
	--------------
	signal RX_L_3, TX_L_3:  std_logic_vector (31 downto 0);
	signal RTS_L_3, DRTS_L_3, CTS_L_3, DCTS_L_3: std_logic;
	--------------
	signal RX_L_4, TX_L_4:  std_logic_vector (31 downto 0);
	signal RTS_L_4, DRTS_L_4, CTS_L_4, DCTS_L_4: std_logic;
	--------------
	signal RX_L_5, TX_L_5:  std_logic_vector (31 downto 0);
	signal RTS_L_5, DRTS_L_5, CTS_L_5, DCTS_L_5: std_logic;
	--------------
	signal RX_L_6, TX_L_6:  std_logic_vector (31 downto 0);
	signal RTS_L_6, DRTS_L_6, CTS_L_6, DCTS_L_6: std_logic;
	--------------
	signal RX_L_7, TX_L_7:  std_logic_vector (31 downto 0);
	signal RTS_L_7, DRTS_L_7, CTS_L_7, DCTS_L_7: std_logic;
	--------------
	signal RX_L_8, TX_L_8:  std_logic_vector (31 downto 0);
	signal RTS_L_8, DRTS_L_8, CTS_L_8, DCTS_L_8: std_logic;
	--------------
	signal RX_L_9, TX_L_9:  std_logic_vector (31 downto 0);
	signal RTS_L_9, DRTS_L_9, CTS_L_9, DCTS_L_9: std_logic;
	--------------
	signal RX_L_10, TX_L_10:  std_logic_vector (31 downto 0);
	signal RTS_L_10, DRTS_L_10, CTS_L_10, DCTS_L_10: std_logic;
	--------------
	signal RX_L_11, TX_L_11:  std_logic_vector (31 downto 0);
	signal RTS_L_11, DRTS_L_11, CTS_L_11, DCTS_L_11: std_logic;
	--------------
	signal RX_L_12, TX_L_12:  std_logic_vector (31 downto 0);
	signal RTS_L_12, DRTS_L_12, CTS_L_12, DCTS_L_12: std_logic;
	--------------
	signal RX_L_13, TX_L_13:  std_logic_vector (31 downto 0);
	signal RTS_L_13, DRTS_L_13, CTS_L_13, DCTS_L_13: std_logic;
	--------------
	signal RX_L_14, TX_L_14:  std_logic_vector (31 downto 0);
	signal RTS_L_14, DRTS_L_14, CTS_L_14, DCTS_L_14: std_logic;
	--------------
	signal RX_L_15, TX_L_15:  std_logic_vector (31 downto 0);
	signal RTS_L_15, DRTS_L_15, CTS_L_15, DCTS_L_15: std_logic;
	--------------
 constant clk_period : time := 1 ns;
signal reset,clk: std_logic :='0';

begin

   clk_process :process
   begin
        clk <= '0';
        wait for clk_period/2;   
        clk <= '1';
        wait for clk_period/2; 
   end process;

reset <= '1' after 1 ns;
-- instantiating the network
NoC: network_4x4 generic map (DATA_WIDTH  => 32)
PORT MAP (reset, clk, 
	RX_L_0, RTS_L_0, CTS_L_0, DRTS_L_0, DCTS_L_0, TX_L_0,
	RX_L_1, RTS_L_1, CTS_L_1, DRTS_L_1, DCTS_L_1, TX_L_1,
	RX_L_2, RTS_L_2, CTS_L_2, DRTS_L_2, DCTS_L_2, TX_L_2,
	RX_L_3, RTS_L_3, CTS_L_3, DRTS_L_3, DCTS_L_3, TX_L_3,
	RX_L_4, RTS_L_4, CTS_L_4, DRTS_L_4, DCTS_L_4, TX_L_4,
	RX_L_5, RTS_L_5, CTS_L_5, DRTS_L_5, DCTS_L_5, TX_L_5,
	RX_L_6, RTS_L_6, CTS_L_6, DRTS_L_6, DCTS_L_6, TX_L_6,
	RX_L_7, RTS_L_7, CTS_L_7, DRTS_L_7, DCTS_L_7, TX_L_7,
	RX_L_8, RTS_L_8, CTS_L_8, DRTS_L_8, DCTS_L_8, TX_L_8,
	RX_L_9, RTS_L_9, CTS_L_9, DRTS_L_9, DCTS_L_9, TX_L_9,
	RX_L_10, RTS_L_10, CTS_L_10, DRTS_L_10, DCTS_L_10, TX_L_10,
	RX_L_11, RTS_L_11, CTS_L_11, DRTS_L_11, DCTS_L_11, TX_L_11,
	RX_L_12, RTS_L_12, CTS_L_12, DRTS_L_12, DCTS_L_12, TX_L_12,
	RX_L_13, RTS_L_13, CTS_L_13, DRTS_L_13, DCTS_L_13, TX_L_13,
	RX_L_14, RTS_L_14, CTS_L_14, DRTS_L_14, DCTS_L_14, TX_L_14,
	RX_L_15, RTS_L_15, CTS_L_15, DRTS_L_15, DCTS_L_15, TX_L_15);

-- connecting the packet generators
gen_packet(9, 0, 10, 1, 2, clk, CTS_L_0, DRTS_L_0, RX_L_0);
gen_packet(6, 1, 12, 1, 2, clk, CTS_L_1, DRTS_L_1, RX_L_1);
gen_packet(8, 2, 11, 1, 2, clk, CTS_L_2, DRTS_L_2, RX_L_2);
gen_packet(4, 3, 10, 1, 2, clk, CTS_L_3, DRTS_L_3, RX_L_3);
gen_packet(10, 4, 3, 1, 2, clk, CTS_L_4, DRTS_L_4, RX_L_4);
gen_packet(7, 5, 9, 1, 2, clk, CTS_L_5, DRTS_L_5, RX_L_5);
gen_packet(10, 6, 1, 1, 2, clk, CTS_L_6, DRTS_L_6, RX_L_6);
gen_packet(5, 7, 13, 1, 2, clk, CTS_L_7, DRTS_L_7, RX_L_7);
gen_packet(4, 8, 11, 1, 2, clk, CTS_L_8, DRTS_L_8, RX_L_8);
gen_packet(4, 9, 12, 1, 2, clk, CTS_L_9, DRTS_L_9, RX_L_9);
gen_packet(3, 10, 11, 1, 2, clk, CTS_L_10, DRTS_L_10, RX_L_10);
gen_packet(6, 11, 4, 1, 2, clk, CTS_L_11, DRTS_L_11, RX_L_11);
gen_packet(4, 12, 6, 1, 2, clk, CTS_L_12, DRTS_L_12, RX_L_12);
gen_packet(10, 13, 6, 1, 2, clk, CTS_L_13, DRTS_L_13, RX_L_13);
gen_packet(6, 14, 0, 1, 2, clk, CTS_L_14, DRTS_L_14, RX_L_14);
gen_packet(9, 15, 8, 1, 2, clk, CTS_L_15, DRTS_L_15, RX_L_15);

-- connecting the packet receivers
get_packet(32, 5,  clk, DCTS_L_0, RTS_L_0, TX_L_0);
get_packet(32, 5,  clk, DCTS_L_1, RTS_L_1, TX_L_1);
get_packet(32, 5,  clk, DCTS_L_2, RTS_L_2, TX_L_2);
get_packet(32, 5,  clk, DCTS_L_3, RTS_L_3, TX_L_3);
get_packet(32, 5,  clk, DCTS_L_4, RTS_L_4, TX_L_4);
get_packet(32, 5,  clk, DCTS_L_5, RTS_L_5, TX_L_5);
get_packet(32, 5,  clk, DCTS_L_6, RTS_L_6, TX_L_6);
get_packet(32, 5,  clk, DCTS_L_7, RTS_L_7, TX_L_7);
get_packet(32, 5,  clk, DCTS_L_8, RTS_L_8, TX_L_8);
get_packet(32, 5,  clk, DCTS_L_9, RTS_L_9, TX_L_9);
get_packet(32, 5,  clk, DCTS_L_10, RTS_L_10, TX_L_10);
get_packet(32, 5,  clk, DCTS_L_11, RTS_L_11, TX_L_11);
get_packet(32, 5,  clk, DCTS_L_12, RTS_L_12, TX_L_12);
get_packet(32, 5,  clk, DCTS_L_13, RTS_L_13, TX_L_13);
get_packet(32, 5,  clk, DCTS_L_14, RTS_L_14, TX_L_14);
get_packet(32, 5,  clk, DCTS_L_15, RTS_L_15, TX_L_15);
end;

