--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated!
-- Here are the parameters:
-- 	 network size x: 2
-- 	 network size y: 2
-- 	 Data width: 32
-- 	 Parity: False
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.numeric_std.ALL;
use work.component_pack.all;

entity network_2x2_with_PE is
 generic (DATA_WIDTH: integer := 32;
          DATA_WIDTH_LV: integer := 11;
          memory_type : string :=
            "TRI_PORT_X"
           --   "DUAL_PORT_"
           --   "ALTERA_LPM"
           --   "XILINX_16X"
      );

port (reset: in  std_logic;
      clk: in  std_logic;

      -- IJTAG network for fault injection and checker status monitoring
      TCK         : in std_logic;
      RST         : in std_logic;
      SEL         : in std_logic;
      SI          : in std_logic;
      SE          : in std_logic;
      UE          : in std_logic;
      CE          : in std_logic;
      SO          : out std_logic;
      toF         : out std_logic;
      toC         : out std_logic;

      -- GPIO for Node 0
      GPIO_out: out  std_logic_vector(15 downto 0);
      GPIO_in: in  std_logic_vector(21 downto 0);

      -- UART for all Plasmas
      uart_write_0  : out std_logic;
      uart_read_0   : in std_logic;
      uart_write_1  : out std_logic;
      uart_read_1   : in std_logic;
      uart_write_2  : out std_logic;
      uart_read_2   : in std_logic;
      uart_write_3  : out std_logic;
      uart_read_3   : in std_logic;

      -- Monitor connections
      temperature_control   : out std_logic_vector(2 downto 0);
      iddt_control          : out std_logic_vector(2 downto 0);
      slack_control         : out std_logic_vector(2 downto 0);
      slack_data            : in std_logic_vector(31 downto 0);
      voltage_control       : out std_logic_vector(2 downto 0);
      voltage_data          : in std_logic_vector(31 downto 0)
    );

end network_2x2_with_PE;


architecture behavior of network_2x2_with_PE is

constant RAMDataSize : positive := 32;
constant RAMAddrSize : positive := 12;
constant path : string(1 to 12) := "Testbenches/"; --uncomment this if you are SIMULATING in MODELSIM, or if you're synthesizing.
-- constant path : string(positive range <>) := "/home/tsotne/ownCloud/git/Bonfire_sim/Bonfire/RTL/Chip_Designs/IMMORTAL_Chip_2017/Testbenches/"; --used only for Vivado similation. Tsotnes PC.

component immortal_sensor_IJTAG_interface is
    Port ( -- Scan Interface  client --------------
            TCK         : in std_logic;
            RST         : in std_logic;
            SEL         : in std_logic;
            SI          : in std_logic;
            SE          : in std_logic;
            UE          : in std_logic;
            CE          : in std_logic;
            SO          : out std_logic;
            toF         : out std_logic;
            toC         : out std_logic;

            -- Monitor connections
            temperature_control   : out std_logic_vector(2 downto 0);
            temperature_data      : in std_logic_vector(12 downto 0);
            iddt_control          : out std_logic_vector(2 downto 0);
            iddt_data             : in std_logic_vector(12 downto 0);
            slack_control         : out std_logic_vector(2 downto 0);
            slack_data            : in std_logic_vector(31 downto 0);
            voltage_control       : out std_logic_vector(2 downto 0);
            voltage_data          : in std_logic_vector(31 downto 0));
end component;

component SIB_mux_pre_FCX_SELgate is
    Port ( -- Scan Interface  client --------------
           SI : in STD_LOGIC; -- ScanInPort
           CE : in STD_LOGIC; -- CaptureEnPort
           SE : in STD_LOGIC; -- ShiftEnPort
           UE : in STD_LOGIC; -- UpdateEnPort
           SEL : in STD_LOGIC; -- SelectPort
           RST : in STD_LOGIC; -- ResetPort
           TCK : in STD_LOGIC; -- TCKPort
           SO : out STD_LOGIC; -- ScanOutPort
           toF : out STD_LOGIC; -- To F flag of the upper hierarchical level
           toC : out STD_LOGIC; -- To C flag of the upper hierarchical level
       -- Scan Interface  host ----------------
           fromSO : in  STD_LOGIC; -- ScanInPort
           toCE : out  STD_LOGIC; -- ToCaptureEnPort
           toSE : out  STD_LOGIC; -- ToShiftEnPort
           toUE : out  STD_LOGIC; -- ToUpdateEnPort
           toSEL : out  STD_LOGIC; -- ToSelectPort
           toRST : out  STD_LOGIC; -- ToResetPort
           toTCK : out  STD_LOGIC; -- ToTCKPort
           toSI : out  STD_LOGIC; -- ScanOutPort
           fromF : in STD_LOGIC; -- From an OR of all F flags in the underlying network segment
           fromC : in STD_LOGIC);  -- From an AND of all C flags in the underlying network segment
end component;

component RAMAccessInstrument is
    Generic ( DataSize : positive := 8;
            AddressSize : positive := 8);
    Port ( -- Scan Interface scan_client ----------
            SI : in std_logic; -- ScanInPort
            SO : out std_logic; -- ScanOutPort
            SEL : in std_logic; -- SelectPort
            ----------------------------------------
            SE : in std_logic; -- ShiftEnPort
            CE : in std_logic; -- CaptureEnPort
            UE : in std_logic; -- UpdateEnPort
            RST : in std_logic; -- ResetPort
            TCK : in std_logic; -- TCKPort
            MEM_SIB_SEL : out std_logic;
               -- RAM interface
            RAM_data_read : in std_logic_vector (DataSize-1 downto 0);
            RAM_data_write : out std_logic_vector (DataSize-1 downto 0);
            RAM_address_out : out std_logic_vector (AddressSize-1 downto 0);
            RAM_write_enable : out std_logic);
end component;

-- Monitor signals
signal temperature_data      : std_logic_vector(12 downto 0);
signal iddt_data             : std_logic_vector(12 downto 0);


-- Declaring network component

-- Declaring NoC_Node component (with Plasma, RAM, NI and UART)


-- generating bulk signals...
    signal RX_L_0, TX_L_0:  std_logic_vector (31 downto 0);
    signal credit_counter_out_0:  std_logic_vector (1 downto 0);
    signal credit_out_L_0, credit_in_L_0, valid_in_L_0, valid_out_L_0: std_logic;
    signal RX_L_1, TX_L_1:  std_logic_vector (31 downto 0);
    signal credit_counter_out_1:  std_logic_vector (1 downto 0);
    signal credit_out_L_1, credit_in_L_1, valid_in_L_1, valid_out_L_1: std_logic;
    signal RX_L_2, TX_L_2:  std_logic_vector (31 downto 0);
    signal credit_counter_out_2:  std_logic_vector (1 downto 0);
    signal credit_out_L_2, credit_in_L_2, valid_in_L_2, valid_out_L_2: std_logic;
    signal RX_L_3, TX_L_3:  std_logic_vector (31 downto 0);
    signal credit_counter_out_3:  std_logic_vector (1 downto 0);
    signal credit_out_L_3, credit_in_L_3, valid_in_L_3, valid_out_L_3: std_logic;

    -- NI testing signals
    --------------
    --signal Rxy_reconf: std_logic_vector (7 downto 0) := "01111101";
    --signal Reconfig: std_logic := '0';
    --------------

    signal not_reset: std_logic;

    signal link_faults_0, link_faults_1, link_faults_2, link_faults_3   : std_logic_vector(4 downto 0);
    signal turn_faults_0, turn_faults_1, turn_faults_2, turn_faults_3   : std_logic_vector(19 downto 0);
    signal Rxy_reconf_PE_0, Rxy_reconf_PE_1,Rxy_reconf_PE_2, Rxy_reconf_PE_3   : std_logic_vector(7 downto 0);
    signal Cx_reconf_PE_0, Cx_reconf_PE_1, Cx_reconf_PE_2, Cx_reconf_PE_3 : std_logic_vector(3 downto 0);
    signal Reconfig_command_0, Reconfig_command_1, Reconfig_command_2, Reconfig_command_3 : std_logic;

    signal GPIO_out_FF_in, GPIO_out_FF : std_logic_vector(15 downto 0);
    signal UART_0_W_in, UART_0_W_out, UART_0_R_in, UART_0_R_out : std_logic;
    signal UART_1_W_in, UART_1_W_out, UART_1_R_in, UART_1_R_out : std_logic;
    signal UART_2_W_in, UART_2_W_out, UART_2_R_in, UART_2_R_out : std_logic;
    signal UART_3_W_in, UART_3_W_out, UART_3_R_in, UART_3_R_out : std_logic;

    -- IJTAG-related signals

    signal SO_NoC , SO_sensors , SO_RAM  : std_logic;
    signal toF_NoC, toF_sensors, toF_RAM : std_logic;
    signal toC_NoC, toC_sensors, toC_RAM : std_logic;

    signal SIB_RAM_toSI, SIB_RAM_toTCK, SIB_RAM_toRST, SIB_RAM_toSEL, SIB_RAM_toUE, SIB_RAM_toSE, SIB_RAM_toCE : std_logic;
    signal RAM0_SO,           RAM1_SO,           RAM2_SO,           RAM3_SO           : std_logic;
    signal RAM0_write_enable, RAM1_write_enable, RAM2_write_enable, RAM3_write_enable : std_logic;
    signal RAM0_address,      RAM1_address,      RAM2_address,      RAM3_address      : std_logic_vector(RAMAddrSize-1 downto 0);

    signal IJTAG_ram_0_select            : std_logic;
    signal IJTAG_ram_0_clk               : std_logic;
    signal IJTAG_ram_0_reset             : std_logic;
    signal IJTAG_ram_0_enable            : std_logic;
    signal IJTAG_ram_0_write_byte_enable : std_logic_vector(3 downto 0);
    signal IJTAG_ram_0_address           : std_logic_vector(31 downto 2);
    signal IJTAG_ram_0_data_write        : std_logic_vector(31 downto 0);
    signal IJTAG_ram_0_data_read         : std_logic_vector(31 downto 0);

    signal IJTAG_ram_1_select            : std_logic;
    signal IJTAG_ram_1_clk               : std_logic;
    signal IJTAG_ram_1_reset             : std_logic;
    signal IJTAG_ram_1_enable            : std_logic;
    signal IJTAG_ram_1_write_byte_enable : std_logic_vector(3 downto 0);
    signal IJTAG_ram_1_address           : std_logic_vector(31 downto 2);
    signal IJTAG_ram_1_data_write        : std_logic_vector(31 downto 0);
    signal IJTAG_ram_1_data_read         : std_logic_vector(31 downto 0);

    signal IJTAG_ram_2_select            : std_logic;
    signal IJTAG_ram_2_clk               : std_logic;
    signal IJTAG_ram_2_reset             : std_logic;
    signal IJTAG_ram_2_enable            : std_logic;
    signal IJTAG_ram_2_write_byte_enable : std_logic_vector(3 downto 0);
    signal IJTAG_ram_2_address           : std_logic_vector(31 downto 2);
    signal IJTAG_ram_2_data_write        : std_logic_vector(31 downto 0);
    signal IJTAG_ram_2_data_read         : std_logic_vector(31 downto 0);

    signal IJTAG_ram_3_select            : std_logic;
    signal IJTAG_ram_3_clk               : std_logic;
    signal IJTAG_ram_3_reset             : std_logic;
    signal IJTAG_ram_3_enable            : std_logic;
    signal IJTAG_ram_3_write_byte_enable : std_logic_vector(3 downto 0);
    signal IJTAG_ram_3_address           : std_logic_vector(31 downto 2);
    signal IJTAG_ram_3_data_write        : std_logic_vector(31 downto 0);
    signal IJTAG_ram_3_data_read         : std_logic_vector(31 downto 0);
begin

-- instantiating the network
NoC: network_2x2 generic map (DATA_WIDTH  => 32, DATA_WIDTH_LV => 11)
port map (reset, clk,
    RX_L_0, credit_out_L_0, valid_out_L_0, credit_in_L_0, valid_in_L_0,  TX_L_0,
    RX_L_1, credit_out_L_1, valid_out_L_1, credit_in_L_1, valid_in_L_1,  TX_L_1,
    RX_L_2, credit_out_L_2, valid_out_L_2, credit_in_L_2, valid_in_L_2,  TX_L_2,
    RX_L_3, credit_out_L_3, valid_out_L_3, credit_in_L_3, valid_in_L_3,  TX_L_3,
    link_faults_0, turn_faults_0, Rxy_reconf_PE_0, Cx_reconf_PE_0, Reconfig_command_0,
    link_faults_1, turn_faults_1, Rxy_reconf_PE_1, Cx_reconf_PE_1, Reconfig_command_1,
    link_faults_2, turn_faults_2, Rxy_reconf_PE_2, Cx_reconf_PE_2, Reconfig_command_2,
    link_faults_3, turn_faults_3, Rxy_reconf_PE_3, Cx_reconf_PE_3, Reconfig_command_3,
    TCK, RST, SEL, SO_sensors, SE, UE, CE, SO_NoC, toF_NoC, toC_NoC
    );

process (not_reset, clk)
begin
  if not_reset = '1' then
      GPIO_out_FF <= (others => '0');

      UART_0_W_out <= '0';
      UART_1_W_out <= '0';
      UART_2_W_out <= '0';
      UART_3_W_out <= '0';

      UART_0_R_out <= '0';
      UART_1_R_out <= '0';
      UART_2_R_out <= '0';
      UART_3_R_out <= '0';

  elsif clk'event and clk = '1' then
      GPIO_out_FF <= GPIO_out_FF_in;

      UART_0_W_out <= UART_0_W_in;
      UART_1_W_out <= UART_1_W_in;
      UART_2_W_out <= UART_2_W_in;
      UART_3_W_out <= UART_3_W_in;

      UART_0_R_out <= UART_0_R_in;
      UART_1_R_out <= UART_1_R_in;
      UART_2_R_out <= UART_2_R_in;
      UART_3_R_out <= UART_3_R_in;
  end if;
end process;


GPIO_out <=  GPIO_out_FF;

uart_write_0 <= UART_0_W_out;
uart_write_1 <= UART_1_W_out;
uart_write_2 <= UART_2_W_out;
uart_write_3 <= UART_3_W_out;

UART_0_R_in <= uart_read_0;
UART_1_R_in <= uart_read_1;
UART_2_R_in <= uart_read_2;
UART_3_R_in <= uart_read_3;

not_reset <= not reset;

-- instantiating and connecting the PEs
PE_0: NoC_Node
generic map( current_address => 0,
    stim_file => path & "code_0.txt",
    log_file  => path & "output_0.txt",
    memory_type => memory_type)

port map( not_reset, clk,
        uart_read         => UART_0_R_out,
        uart_write        => UART_0_W_in,
        credit_in => credit_out_L_0,
        valid_out => valid_in_L_0,
        TX => RX_L_0,

        credit_out => credit_in_L_0,
        valid_in => valid_out_L_0,
        RX => TX_L_0,
        link_faults         => link_faults_0,
        turn_faults         => turn_faults_0,
        Rxy_reconf_PE       => Rxy_reconf_PE_0,
        Cx_reconf_PE        => Cx_reconf_PE_0,
        Reconfig_command    => Reconfig_command_0,

        GPIO_out            => GPIO_out_FF_in,
        GPIO_in             => GPIO_in,
        IJTAG_select            => IJTAG_ram_0_select,
        IJTAG_clk               => IJTAG_ram_0_clk,
        IJTAG_reset             => IJTAG_ram_0_reset,
        IJTAG_enable            => IJTAG_ram_0_enable,
        IJTAG_write_byte_enable => IJTAG_ram_0_write_byte_enable,
        IJTAG_address           => IJTAG_ram_0_address,
        IJTAG_data_write        => IJTAG_ram_0_data_write,
        IJTAG_data_read         => IJTAG_ram_0_data_read
   );

PE_1: NoC_Node
generic map( current_address => 1,
    stim_file => path & "code_1.txt",
    log_file  => path & "output_1.txt",
    memory_type => memory_type)

port map( not_reset, clk,
        uart_read         => UART_1_R_out,
        uart_write        => UART_1_W_in,

        credit_in => credit_out_L_1,
        valid_out => valid_in_L_1,
        TX => RX_L_1,

        credit_out => credit_in_L_1,
        valid_in => valid_out_L_1,
        RX => TX_L_1,
        link_faults         => link_faults_1,
        turn_faults         => turn_faults_1,
        Rxy_reconf_PE       => Rxy_reconf_PE_1,
        Cx_reconf_PE        => Cx_reconf_PE_1,
        Reconfig_command    => Reconfig_command_1,

        GPIO_out            => open,
        GPIO_in             => (others => '0'),

        IJTAG_select            => IJTAG_ram_1_select,
        IJTAG_clk               => IJTAG_ram_1_clk,
        IJTAG_reset             => IJTAG_ram_1_reset,
        IJTAG_enable            => IJTAG_ram_1_enable,
        IJTAG_write_byte_enable => IJTAG_ram_1_write_byte_enable,
        IJTAG_address           => IJTAG_ram_1_address,
        IJTAG_data_write        => IJTAG_ram_1_data_write,
        IJTAG_data_read         => IJTAG_ram_1_data_read
   );

PE_2: NoC_Node
generic map( current_address => 2,
    stim_file => path & "code_2.txt",
    log_file  => path & "output_2.txt",
    memory_type => memory_type)

port map( not_reset, clk,
        uart_read         => UART_2_R_out,
        uart_write        => UART_2_W_in,

        credit_in => credit_out_L_2,
        valid_out => valid_in_L_2,
        TX => RX_L_2,

        credit_out => credit_in_L_2,
        valid_in => valid_out_L_2,
        RX => TX_L_2,
        link_faults         => link_faults_2,
        turn_faults         => turn_faults_2,
        Rxy_reconf_PE       => Rxy_reconf_PE_2,
        Cx_reconf_PE        => Cx_reconf_PE_2,
        Reconfig_command    => Reconfig_command_2,

        GPIO_out            => open,
        GPIO_in             => (others => '0'),
        IJTAG_select            => IJTAG_ram_2_select,
        IJTAG_clk               => IJTAG_ram_2_clk,
        IJTAG_reset             => IJTAG_ram_2_reset,
        IJTAG_enable            => IJTAG_ram_2_enable,
        IJTAG_write_byte_enable => IJTAG_ram_2_write_byte_enable,
        IJTAG_address           => IJTAG_ram_2_address,
        IJTAG_data_write        => IJTAG_ram_2_data_write,
        IJTAG_data_read         => IJTAG_ram_2_data_read
   );

PE_3: NoC_Node
generic map( current_address => 3,
    stim_file => path & "code_3.txt",
    log_file  => path & "output_3.txt",
    memory_type => memory_type)

port map( not_reset, clk,
        uart_read         => UART_3_R_out,
        uart_write        => UART_3_W_in,

        credit_in => credit_out_L_3,
        valid_out => valid_in_L_3,
        TX => RX_L_3,

        credit_out => credit_in_L_3,
        valid_in => valid_out_L_3,
        RX => TX_L_3,
        link_faults         => link_faults_3,
        turn_faults         => turn_faults_3,
        Rxy_reconf_PE       => Rxy_reconf_PE_3,
        Cx_reconf_PE        => Cx_reconf_PE_3,
        Reconfig_command    => Reconfig_command_3,

        GPIO_out            => open,
        GPIO_in             => (others => '0'),
        IJTAG_select            => IJTAG_ram_3_select,
        IJTAG_clk               => IJTAG_ram_3_clk,
        IJTAG_reset             => IJTAG_ram_3_reset,
        IJTAG_enable            => IJTAG_ram_3_enable,
        IJTAG_write_byte_enable => IJTAG_ram_3_write_byte_enable,
        IJTAG_address           => IJTAG_ram_3_address,
        IJTAG_data_write        => IJTAG_ram_3_data_write,
        IJTAG_data_read         => IJTAG_ram_3_data_read
   );

-------------------------------------------
------- IJTAG stuff -----------------------
-------------------------------------------

--   Organization of IJTAG network (top level):
--            .----------.   .-----------.   .----------.
--     SI ----| sib_ram  |---| sib_sens  |---| sib_noc  |-- SO
--            '----------'   '-----------'   '----------'
--              |       |_________________________________________________.
--              |                                                         |
--              | .-----------. .-----------. .-----------. .-----------. |
--              '-| sib_ram_0 |-| sib_ram_1 |-| sib_ram_2 |-| sib_ram_3 |-'
--                '-----------' '-----------' '-----------' '-----------'

toF <= toF_NoC or toF_sensors;
toC <= toC_NoC and toC_sensors;
SO <= SO_NoC;

IJTAG_ram_0_enable <= '1';
IJTAG_ram_1_enable <= '1';
IJTAG_ram_2_enable <= '1';
IJTAG_ram_3_enable <= '1';

IJTAG_ram_0_clk <= TCK;
IJTAG_ram_1_clk <= TCK;
IJTAG_ram_2_clk <= TCK;
IJTAG_ram_3_clk <= TCK;

IJTAG_ram_0_reset <= RST;
IJTAG_ram_1_reset <= RST;
IJTAG_ram_2_reset <= RST;
IJTAG_ram_3_reset <= RST;

-- RAM Access SIB

SIB_RAM : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI  => SI,
    CE  => CE,
    SE  => SE,
    UE  => UE,
    SEL => SEL,
    RST => RST,
    TCK => TCK,
    SO  => SO_RAM,
    toF => toF_RAM,
    toC => toC_RAM,
     -- Scan Interface  host ----------------
    fromSO => RAM3_SO,
    toCE   => SIB_RAM_toCE,
    toSE   => SIB_RAM_toSE,
    toUE   => SIB_RAM_toUE,
    toSEL  => SIB_RAM_toSEL,
    toRST  => SIB_RAM_toRST,
    toTCK  => SIB_RAM_toTCK,
    toSI   => SIB_RAM_toSI,
    fromF  => '0',
    fromC  => '1'
);

-- RAM Access instruments

RAM_instr0 : RAMAccessInstrument
 generic map ( DataSize => RAMDataSize,
               AddressSize => RAMAddrSize)
    port map ( SI  => SIB_RAM_toSI,
               SO  => RAM0_SO,
               SEL => SIB_RAM_toSEL,
               SE  => SIB_RAM_toSE,
               CE  => SIB_RAM_toCE,
               UE  => SIB_RAM_toUE,
               RST => SIB_RAM_toRST,
               TCK => SIB_RAM_toTCK,
               MEM_SIB_SEL => IJTAG_ram_0_select,
               RAM_data_read => IJTAG_ram_0_data_read,
               RAM_data_write => IJTAG_ram_0_data_write,
               RAM_address_out => RAM0_address,
               RAM_write_enable => RAM0_write_enable);

IJTAG_ram_0_write_byte_enable <= (others => RAM0_write_enable);
IJTAG_ram_0_address <= "000000000000000000" & RAM0_address;

RAM_instr1 : RAMAccessInstrument
 generic map ( DataSize => RAMDataSize,
               AddressSize => RAMAddrSize)
    port map ( SI  => RAM0_SO,
               SO  => RAM1_SO,
               SEL => SIB_RAM_toSEL,
               SE  => SIB_RAM_toSE,
               CE  => SIB_RAM_toCE,
               UE  => SIB_RAM_toUE,
               RST => SIB_RAM_toRST,
               TCK => SIB_RAM_toTCK,
               MEM_SIB_SEL => IJTAG_ram_1_select,
               RAM_data_read => IJTAG_ram_1_data_read,
               RAM_data_write => IJTAG_ram_1_data_write,
               RAM_address_out => RAM1_address,
               RAM_write_enable => RAM1_write_enable);

IJTAG_ram_1_write_byte_enable <= (others => RAM1_write_enable);
IJTAG_ram_1_address <= "000000000000000000" & RAM1_address;

RAM_instr2 : RAMAccessInstrument
 generic map ( DataSize => RAMDataSize,
               AddressSize => RAMAddrSize)
    port map ( SI  => RAM1_SO,
               SO  => RAM2_SO,
               SEL => SIB_RAM_toSEL,
               SE  => SIB_RAM_toSE,
               CE  => SIB_RAM_toCE,
               UE  => SIB_RAM_toUE,
               RST => SIB_RAM_toRST,
               TCK => SIB_RAM_toTCK,
               MEM_SIB_SEL => IJTAG_ram_2_select,
               RAM_data_read => IJTAG_ram_2_data_read,
               RAM_data_write => IJTAG_ram_2_data_write,
               RAM_address_out => RAM2_address,
               RAM_write_enable => RAM2_write_enable);

IJTAG_ram_2_write_byte_enable <= (others => RAM2_write_enable);
IJTAG_ram_2_address <= "000000000000000000" & RAM2_address;

RAM_instr3 : RAMAccessInstrument
 generic map ( DataSize => RAMDataSize,
               AddressSize => RAMAddrSize)
    port map ( SI  => RAM2_SO,
               SO  => RAM3_SO,
               SEL => SIB_RAM_toSEL,
               SE  => SIB_RAM_toSE,
               CE  => SIB_RAM_toCE,
               UE  => SIB_RAM_toUE,
               RST => SIB_RAM_toRST,
               TCK => SIB_RAM_toTCK,
               MEM_SIB_SEL => IJTAG_ram_3_select,
               RAM_data_read => IJTAG_ram_3_data_read,
               RAM_data_write => IJTAG_ram_3_data_write,
               RAM_address_out => RAM3_address,
               RAM_write_enable => RAM3_write_enable);

IJTAG_ram_3_write_byte_enable <= (others => RAM3_write_enable);
IJTAG_ram_3_address <= "000000000000000000" & RAM3_address;

-- IMMORTAL sensors interface

immortal_sensors: immortal_sensor_IJTAG_interface
    port map (
    TCK => TCK,
    RST => RST,
    SEL => SEL,
    SI  => SO_RAM,
    SE  => SE,
    UE  => UE,
    CE  => CE,
    SO  => SO_sensors,
    toF => toF_sensors,
    toC => toC_sensors,

    temperature_control => temperature_control,
    temperature_data    => temperature_data,
    iddt_control        => iddt_control,
    iddt_data           => iddt_data,
    slack_control       => slack_control,
    slack_data          => slack_data,
    voltage_control     => voltage_control,
    voltage_data        => voltage_data
  );

temperature_data <= (others => '0');
iddt_data <= (others => '0');

end;
