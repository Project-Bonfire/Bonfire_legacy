--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated!
-- Here are the parameters:
-- 	 network size x: 2
-- 	 network size y: 2
-- 	 Data width: 32
-- 	 Parity: False
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.numeric_std.ALL; 

entity network_2x2 is
 generic (DATA_WIDTH: integer := 32; DATA_WIDTH_LV: integer := 11);
port (reset: in  std_logic; 
	clk: in  std_logic; 
	--------------
	--------------
	RX_L_0: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_0, valid_out_L_0: out std_logic;
	credit_in_L_0, valid_in_L_0: in std_logic;
	TX_L_0: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_1: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_1, valid_out_L_1: out std_logic;
	credit_in_L_1, valid_in_L_1: in std_logic;
	TX_L_1: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_2: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_2, valid_out_L_2: out std_logic;
	credit_in_L_2, valid_in_L_2: in std_logic;
	TX_L_2: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_3: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_3, valid_out_L_3: out std_logic;
	credit_in_L_3, valid_in_L_3: in std_logic;
	TX_L_3: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
    link_faults_0: out std_logic_vector(4 downto 0);
    turn_faults_0: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_0: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_0: in  std_logic_vector(3 downto 0);
    Reconfig_command_0 : in std_logic;

	--------------
    link_faults_1: out std_logic_vector(4 downto 0);
    turn_faults_1: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_1: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_1: in  std_logic_vector(3 downto 0);
    Reconfig_command_1 : in std_logic;

	--------------
    link_faults_2: out std_logic_vector(4 downto 0);
    turn_faults_2: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_2: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_2: in  std_logic_vector(3 downto 0);
    Reconfig_command_2 : in std_logic;

	--------------
    link_faults_3: out std_logic_vector(4 downto 0);
    turn_faults_3: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_3: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_3: in  std_logic_vector(3 downto 0);
    Reconfig_command_3 : in std_logic; 

    --------------
    -- IJTAG network for fault injection and checker status monitoring
    TCK         : in std_logic;
    RST         : in std_logic;
    SEL         : in std_logic;
    SI          : in std_logic;
    SE          : in std_logic;
    UE          : in std_logic;
    CE          : in std_logic;
    SO          : out std_logic;
    toF         : out std_logic;
    toC         : out std_logic
    ); 
end network_2x2; 


architecture behavior of network_2x2 is

COMPONENT router_credit_based_PD_C_SHMU is  --fault classifier plus packet-dropping 
    generic (
        DATA_WIDTH: integer := 32;
        current_address : integer := 0;
        Rxy_rst : integer := 10;
        Cx_rst : integer := 10;
        healthy_counter_threshold : integer := 8;
        faulty_counter_threshold: integer := 2;
        counter_depth: integer := 4;
        NoC_size: integer := 4
    );
    port (
    reset, clk: in std_logic;

    RX_N, RX_E, RX_W, RX_S, RX_L : in std_logic_vector (DATA_WIDTH-1 downto 0); 
    credit_in_N, credit_in_E, credit_in_W, credit_in_S, credit_in_L: in std_logic;
    valid_in_N, valid_in_E, valid_in_W, valid_in_S, valid_in_L : in std_logic;
    valid_out_N, valid_out_E, valid_out_W, valid_out_S, valid_out_L : out std_logic;
    credit_out_N, credit_out_E, credit_out_W, credit_out_S, credit_out_L: out std_logic;
    TX_N, TX_E, TX_W, TX_S, TX_L: out std_logic_vector (DATA_WIDTH-1 downto 0);

    Faulty_N_in, Faulty_E_in, Faulty_W_in, Faulty_S_in: in std_logic;
    Faulty_N_out, Faulty_E_out, Faulty_W_out, Faulty_S_out: out std_logic;

    -- should be connected to NI
    link_faults: out std_logic_vector(4 downto 0);
    turn_faults: out std_logic_vector(19 downto 0);

    Rxy_reconf_PE: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE: in  std_logic_vector(3 downto 0);
    Reconfig_command : in std_logic;

    -- fault injector shift register with serial input signals
    TCK: in std_logic;  
    SE: in std_logic;       -- shift enable 
    UE: in std_logic;       -- update enable
    SI: in std_logic;       -- serial Input
    SO: out std_logic;      -- serial output

    ---- Outputs for non-classified fault information
    link_faults_async: out std_logic_vector(4 downto 0);
    turn_faults_async: out std_logic_vector(19 downto 0)
 ); 
end COMPONENT; 


-- For IJAG

component SIB_mux_pre_FCX_SELgate is
    Port ( -- Scan Interface  client --------------
           SI : in STD_LOGIC; -- ScanInPort 
           CE : in STD_LOGIC; -- CaptureEnPort
           SE : in STD_LOGIC; -- ShiftEnPort
           UE : in STD_LOGIC; -- UpdateEnPort
           SEL : in STD_LOGIC; -- SelectPort
           RST : in STD_LOGIC; -- ResetPort
           TCK : in STD_LOGIC; -- TCKPort
           SO : out STD_LOGIC; -- ScanOutPort
           toF : out STD_LOGIC; -- To F flag of the upper hierarchical level
           toC : out STD_LOGIC; -- To C flag of the upper hierarchical level
       -- Scan Interface  host ----------------
           fromSO : in  STD_LOGIC; -- ScanInPort
           toCE : out  STD_LOGIC; -- ToCaptureEnPort
           toSE : out  STD_LOGIC; -- ToShiftEnPort
           toUE : out  STD_LOGIC; -- ToUpdateEnPort
           toSEL : out  STD_LOGIC; -- ToSelectPort
           toRST : out  STD_LOGIC; -- ToResetPort
           toTCK : out  STD_LOGIC; -- ToTCKPort
           toSI : out  STD_LOGIC; -- ScanOutPort
           fromF : in STD_LOGIC; -- From an OR of all F flags in the underlying network segment
           fromC : in STD_LOGIC);  -- From an AND of all C flags in the underlying network segment
end component;


-- generating bulk signals. not all of them are used in the design...
	signal credit_out_N_0, credit_out_E_0, credit_out_W_0, credit_out_S_0: std_logic;
	signal credit_out_N_1, credit_out_E_1, credit_out_W_1, credit_out_S_1: std_logic;
	signal credit_out_N_2, credit_out_E_2, credit_out_W_2, credit_out_S_2: std_logic;
	signal credit_out_N_3, credit_out_E_3, credit_out_W_3, credit_out_S_3: std_logic;

	signal credit_in_N_0, credit_in_E_0, credit_in_W_0, credit_in_S_0: std_logic;
	signal credit_in_N_1, credit_in_E_1, credit_in_W_1, credit_in_S_1: std_logic;
	signal credit_in_N_2, credit_in_E_2, credit_in_W_2, credit_in_S_2: std_logic;
	signal credit_in_N_3, credit_in_E_3, credit_in_W_3, credit_in_S_3: std_logic;

	signal RX_N_0, RX_E_0, RX_W_0, RX_S_0 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_1, RX_E_1, RX_W_1, RX_S_1 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_2, RX_E_2, RX_W_2, RX_S_2 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_3, RX_E_3, RX_W_3, RX_S_3 : std_logic_vector (DATA_WIDTH-1 downto 0);

	signal valid_out_N_0, valid_out_E_0, valid_out_W_0, valid_out_S_0: std_logic;
	signal valid_out_N_1, valid_out_E_1, valid_out_W_1, valid_out_S_1: std_logic;
	signal valid_out_N_2, valid_out_E_2, valid_out_W_2, valid_out_S_2: std_logic;
	signal valid_out_N_3, valid_out_E_3, valid_out_W_3, valid_out_S_3: std_logic;

	signal valid_in_N_0, valid_in_E_0, valid_in_W_0, valid_in_S_0: std_logic;
	signal valid_in_N_1, valid_in_E_1, valid_in_W_1, valid_in_S_1: std_logic;
	signal valid_in_N_2, valid_in_E_2, valid_in_W_2, valid_in_S_2: std_logic;
	signal valid_in_N_3, valid_in_E_3, valid_in_W_3, valid_in_S_3: std_logic;

	signal TX_N_0, TX_E_0, TX_W_0, TX_S_0 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_1, TX_E_1, TX_W_1, TX_S_1 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_2, TX_E_2, TX_W_2, TX_S_2 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_3, TX_E_3, TX_W_3, TX_S_3 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal Faulty_N_out0,Faulty_E_out0,Faulty_W_out0,Faulty_S_out0: std_logic;
	signal Faulty_N_in0,Faulty_E_in0,Faulty_W_in0,Faulty_S_in0: std_logic;
	signal Faulty_N_out1,Faulty_E_out1,Faulty_W_out1,Faulty_S_out1: std_logic;
	signal Faulty_N_in1,Faulty_E_in1,Faulty_W_in1,Faulty_S_in1: std_logic;
	signal Faulty_N_out2,Faulty_E_out2,Faulty_W_out2,Faulty_S_out2: std_logic;
	signal Faulty_N_in2,Faulty_E_in2,Faulty_W_in2,Faulty_S_in2: std_logic;
	signal Faulty_N_out3,Faulty_E_out3,Faulty_W_out3,Faulty_S_out3: std_logic;
	signal Faulty_N_in3,Faulty_E_in3,Faulty_W_in3,Faulty_S_in3: std_logic;

    -- fault injector signals
    signal TCK_0, TCK_1, TCK_2, TCK_3: std_logic;
    signal SE_0,  SE_1,  SE_2,  SE_3:  std_logic;
    signal UE_0,  UE_1,  UE_2,  UE_3:  std_logic;
    signal SI_0,  SI_1,  SI_2,  SI_3:  std_logic;
    signal SO_0,  SO_1,  SO_2,  SO_3:  std_logic;

    --------------
    -- IJTAG network signals
    signal SIB_0_toSEL, SIB_1_toSEL, SIB_2_toSEL, SIB_3_toSEL : std_logic;
    signal SIB_0_toCE,  SIB_1_toCE,  SIB_2_toCE,  SIB_3_toCE  : std_logic;
    signal SIB_0_toRST, SIB_1_toRST, SIB_2_toRST, SIB_3_toRST : std_logic;
    signal SIB_0_so,    SIB_1_so,    SIB_2_so,    SIB_3_so    : std_logic;
    -- flags from checkers
    signal F_R0, F_R1, F_R2, F_R3 : std_logic := '0';
    signal C_R0, C_R1, C_R2, C_R3 : std_logic := '1';
    -- flags top level
    signal F_segtop_fromSIB_0, C_segtop_fromSIB_0 : std_logic;
    signal F_segtop_fromSIB_1, C_segtop_fromSIB_1 : std_logic;
    signal F_segtop_fromSIB_2, C_segtop_fromSIB_2 : std_logic;
    signal F_segtop_fromSIB_3, C_segtop_fromSIB_3 : std_logic;
    --------------

    -- the checker output related ports (for unclassified fault information)
    signal link_faults_async_0 : std_logic_vector(4 downto 0);
    signal turn_faults_async_0: std_logic_vector(19 downto 0);

    --------------
    signal link_faults_async_1 : std_logic_vector(4 downto 0);
    signal turn_faults_async_1: std_logic_vector(19 downto 0);

    --------------
    signal link_faults_async_2 : std_logic_vector(4 downto 0);
    signal turn_faults_async_2: std_logic_vector(19 downto 0);

    --------------
    signal link_faults_async_3 : std_logic_vector(4 downto 0);
    signal turn_faults_async_3: std_logic_vector(19 downto 0);
    --------------

    -- Fault injection related signals and constants
    constant fault_clk_period : time := 1 ns;


--        organizaiton of the network:
--     x --------------->
--  y         ----       ----
--  |        | 0  | --- | 1  |
--  |         ----       ----
--  |          |          |
--  |         ----       ----
--  |        | 2  | --- | 3  |
--  v         ----       ----
--                         
begin

   ---- Fault injection clock process (IJTAG-related)
   --fault_clk_process :process
   --begin
   --     TCK_0 <= '0';
   --     wait for fault_clk_period/2;   
   --     TCK_0 <= '1';
   --     wait for fault_clk_period/2; 
   --end process;

   ---- Fault Injection Stimulus process (shifting in single SA0 fault at a location in L FIFO in Router 0)
   --fault_injection_stim_proc: process
   --begin        
   --   wait for 3000 ns;

   --   UE_0 <= '0';
   --   SE_0 <= '1';

   --   -- Not Injecting fault to Allocator logic
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to S Arbiter_out
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to W Arbiter_out
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to E Arbiter_out
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to N Arbiter_out
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to L Arbiter_out
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to S Arbiter_in
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to W Arbiter_in
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to E Arbiter_in
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to N Arbiter_in
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to L Arbiter_in
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to S LBDR
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to W LBDR
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to E LBDR
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to N LBDR
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to L LBDR
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to S FIFO
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA0 fault injection at bit 40 (read_pointer(0))
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA0 fault injection at bit 40 (read_pointer(0))

   --   -- Not Injecting fault to W FIFO
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA1 fault injection at bit 0 (LSB)

   --   -- Injecting fault to E FIFO
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA1 fault injection at bit 0 (LSB)

   --   -- Not Injecting fault to N FIFO
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA1 fault injection at bit 0 (LSB)

   --   -- Injecting fault to L FIFO
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '0'; -- SA1 fault injection at bit 0 (LSB)
   --   wait until TCK_0'event and TCK_0 ='0';
   --     SI_0 <= '1'; -- SA1 fault injection at bit 0 (LSB)

   --   wait until TCK_0'event and TCK_0 ='0'; -- Actually affect the signal(s) with fault information
   --     UE_0 <= '1';
   --     SE_0 <= '0';
   --     SI_0 <= '0'; 
   --   --wait until TCK_0'event and TCK_0 ='0'; -- No fault injection anymore and no shifting

   --   --wait until TCK_0'event and TCK_0 ='0'; -- No fault injection anymore and no shifting
   --   --wait until TCK_0'event and TCK_0 ='0'; -- No fault injection anymore and no shifting
   --   --wait until TCK_0'event and TCK_0 ='0'; -- No fault injection anymore and no shifting
   --   --wait until TCK_0'event and TCK_0 ='0'; -- No fault injection anymore and no shifting
   --   --wait until TCK_0'event and TCK_0 ='0'; -- No fault injection anymore and no shifting

   --   wait until TCK_0'event and TCK_0 ='0'; -- No fault injection anymore and no shifting
   --     UE_0 <= '0';
   --     SE_0 <= '0';
   --     SI_0 <= '0';         
   --   --wait until TCK_0'event and TCK_0 ='0'; 

   --   wait; --??

   --end process;

-- flags top level
toF <= F_segtop_fromSIB_0 or  F_segtop_fromSIB_1 or  F_segtop_fromSIB_2 or  F_segtop_fromSIB_3;
toC <= C_segtop_fromSIB_0 and C_segtop_fromSIB_1 and C_segtop_fromSIB_2 and C_segtop_fromSIB_3;
SO <= SIB_3_so;

SIB_0 : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SI,
    CE => CE,
    SE => SE,
    UE => UE,
    SEL => SEL,
    RST => RST,
    TCK => TCK,
    SO => SIB_0_so,
    toF => F_segtop_fromSIB_0,
    toC => C_segtop_fromSIB_0,
     -- Scan Interface  host ----------------
    fromSO => SO_0,
    toCE => SIB_0_toCE,
    toSE => SE_0,
    toUE => UE_0,
    toSEL => SIB_0_toSEL,
    toRST => SIB_0_toRST,
    toTCK => TCK_0,
    toSI => SI_0,
    fromF => F_R0,
    fromC => C_R0
);
SIB_1 : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_0_so,
    CE => CE,
    SE => SE,
    UE => UE,
    SEL => SEL,
    RST => RST,
    TCK => TCK,
    SO => SIB_1_so,
    toF => F_segtop_fromSIB_1,
    toC => C_segtop_fromSIB_1,
     -- Scan Interface  host ----------------
    fromSO => SO_1,
    toCE => SIB_1_toCE,
    toSE => SE_1,
    toUE => UE_1,
    toSEL => SIB_1_toSEL,
    toRST => SIB_1_toRST,
    toTCK => TCK_1,
    toSI => SI_1,
    fromF => F_R1,
    fromC => C_R1
);
SIB_2 : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_1_so,
    CE => CE,
    SE => SE,
    UE => UE,
    SEL => SEL,
    RST => RST,
    TCK => TCK,
    SO => SIB_2_so,
    toF => F_segtop_fromSIB_2,
    toC => C_segtop_fromSIB_2,
     -- Scan Interface  host ----------------
    fromSO => SO_2,
    toCE => SIB_2_toCE,
    toSE => SE_2,
    toUE => UE_2,
    toSEL => SIB_2_toSEL,
    toRST => SIB_2_toRST,
    toTCK => TCK_2,
    toSI => SI_2,
    fromF => F_R2,
    fromC => C_R2
);
SIB_3 : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_2_so,
    CE => CE,
    SE => SE,
    UE => UE,
    SEL => SEL,
    RST => RST,
    TCK => TCK,
    SO => SIB_3_so,
    toF => F_segtop_fromSIB_3,
    toC => C_segtop_fromSIB_3,
     -- Scan Interface  host ----------------
    fromSO => SO_3,
    toCE => SIB_3_toCE,
    toSE => SE_3,
    toUE => UE_3,
    toSEL => SIB_3_toSEL,
    toRST => SIB_3_toRST,
    toTCK => TCK_3,
    toSI => SI_3,
    fromF => F_R3,
    fromC => C_R3
);


R_0: router_credit_based_PD_C_SHMU 
    generic map (DATA_WIDTH =>DATA_WIDTH,         current_address => 0, Rxy_rst => 60,
        Cx_rst =>  10, NoC_size => 2, healthy_counter_threshold => 15, faulty_counter_threshold => 3, counter_depth => 4)
    port map(
    reset, clk,
	RX_N_0, RX_E_0, RX_W_0, RX_S_0, RX_L_0,
	credit_in_N_0, credit_in_E_0, credit_in_W_0, credit_in_S_0, credit_in_L_0,
	valid_in_N_0, valid_in_E_0, valid_in_W_0, valid_in_S_0, valid_in_L_0,
	valid_out_N_0, valid_out_E_0, valid_out_W_0, valid_out_S_0, valid_out_L_0,
	credit_out_N_0, credit_out_E_0, credit_out_W_0, credit_out_S_0, credit_out_L_0,
	TX_N_0, TX_E_0, TX_W_0, TX_S_0, TX_L_0,
	Faulty_N_in0,Faulty_E_in0,Faulty_W_in0,Faulty_S_in0,
	Faulty_N_out0,Faulty_E_out0,Faulty_W_out0,Faulty_S_out0,
	-- should be connected to NI
	link_faults_0, turn_faults_0,
	Rxy_reconf_PE_0, Cx_reconf_PE_0, Reconfig_command_0, 
	-- fault injector shift register with serial input signals
	TCK_0, SE_0, UE_0, SI_0, SO_0, 
    -- the non-classified fault information
    link_faults_async_0, turn_faults_async_0
 ); 

R_1: router_credit_based_PD_C_SHMU 
    generic map (DATA_WIDTH =>DATA_WIDTH,         current_address => 1, Rxy_rst => 60,
        Cx_rst =>  12, NoC_size => 2, healthy_counter_threshold => 15, faulty_counter_threshold => 3, counter_depth => 4)
    port map(
    reset, clk,
	RX_N_1, RX_E_1, RX_W_1, RX_S_1, RX_L_1,
	credit_in_N_1, credit_in_E_1, credit_in_W_1, credit_in_S_1, credit_in_L_1,
	valid_in_N_1, valid_in_E_1, valid_in_W_1, valid_in_S_1, valid_in_L_1,
	valid_out_N_1, valid_out_E_1, valid_out_W_1, valid_out_S_1, valid_out_L_1,
	credit_out_N_1, credit_out_E_1, credit_out_W_1, credit_out_S_1, credit_out_L_1,
	TX_N_1, TX_E_1, TX_W_1, TX_S_1, TX_L_1,
	Faulty_N_in1,Faulty_E_in1,Faulty_W_in1,Faulty_S_in1,
	Faulty_N_out1,Faulty_E_out1,Faulty_W_out1,Faulty_S_out1,
	-- should be connected to NI
	link_faults_1, turn_faults_1,
	Rxy_reconf_PE_1, Cx_reconf_PE_1, Reconfig_command_1, 
    -- fault injector shift register with serial input signals
    TCK_1, SE_1, UE_1, SI_1, SO_1, 
    -- the non-classified fault information
    link_faults_async_1, turn_faults_async_1
 ); 
R_2: router_credit_based_PD_C_SHMU 
    generic map (DATA_WIDTH =>DATA_WIDTH,         current_address => 2, Rxy_rst => 60,
        Cx_rst =>  3, NoC_size => 2, healthy_counter_threshold => 15, faulty_counter_threshold => 3, counter_depth => 4)
    port map(
    reset, clk,
	RX_N_2, RX_E_2, RX_W_2, RX_S_2, RX_L_2,
	credit_in_N_2, credit_in_E_2, credit_in_W_2, credit_in_S_2, credit_in_L_2,
	valid_in_N_2, valid_in_E_2, valid_in_W_2, valid_in_S_2, valid_in_L_2,
	valid_out_N_2, valid_out_E_2, valid_out_W_2, valid_out_S_2, valid_out_L_2,
	credit_out_N_2, credit_out_E_2, credit_out_W_2, credit_out_S_2, credit_out_L_2,
	TX_N_2, TX_E_2, TX_W_2, TX_S_2, TX_L_2,
	Faulty_N_in2,Faulty_E_in2,Faulty_W_in2,Faulty_S_in2,
	Faulty_N_out2,Faulty_E_out2,Faulty_W_out2,Faulty_S_out2,
	-- should be connected to NI
	link_faults_2, turn_faults_2,
	Rxy_reconf_PE_2, Cx_reconf_PE_2, Reconfig_command_2, 
    -- fault injector shift register with serial input signals
    TCK_2, SE_2, UE_2, SI_2, SO_2, 
    -- the non-classified fault information
    link_faults_async_2, turn_faults_async_2
 ); 
R_3: router_credit_based_PD_C_SHMU 
    generic map (DATA_WIDTH =>DATA_WIDTH,         current_address => 3, Rxy_rst => 60,
        Cx_rst =>  5, NoC_size => 2, healthy_counter_threshold => 15, faulty_counter_threshold => 3, counter_depth => 4)
    port map(
    reset, clk,
	RX_N_3, RX_E_3, RX_W_3, RX_S_3, RX_L_3,
	credit_in_N_3, credit_in_E_3, credit_in_W_3, credit_in_S_3, credit_in_L_3,
	valid_in_N_3, valid_in_E_3, valid_in_W_3, valid_in_S_3, valid_in_L_3,
	valid_out_N_3, valid_out_E_3, valid_out_W_3, valid_out_S_3, valid_out_L_3,
	credit_out_N_3, credit_out_E_3, credit_out_W_3, credit_out_S_3, credit_out_L_3,
	TX_N_3, TX_E_3, TX_W_3, TX_S_3, TX_L_3,
	Faulty_N_in3,Faulty_E_in3,Faulty_W_in3,Faulty_S_in3,
	Faulty_N_out3,Faulty_E_out3,Faulty_W_out3,Faulty_S_out3,
	-- should be connected to NI
	link_faults_3, turn_faults_3,
	Rxy_reconf_PE_3, Cx_reconf_PE_3, Reconfig_command_3, 
    -- fault injector shift register with serial input signals
    TCK_3, SE_3, UE_3, SI_3, SO_3, 
    -- the non-classified fault information
    link_faults_async_3, turn_faults_async_3
 ); 

---------------------------------------------------------------
-- binding the routers together
-- vertical ins/outs
-- connecting router: 0 to router: 2 and vice versa
RX_N_2<= TX_S_0;
RX_S_0<= TX_N_2;
-------------------
-- connecting router: 1 to router: 3 and vice versa
RX_N_3<= TX_S_1;
RX_S_1<= TX_N_3;
-------------------

-- horizontal ins/outs
-- connecting router: 0 to router: 1 and vice versa
RX_E_0 <= TX_W_1;
RX_W_1 <= TX_E_0;
-------------------
-- connecting router: 2 to router: 3 and vice versa
RX_E_2 <= TX_W_3;
RX_W_3 <= TX_E_2;
-------------------
---------------------------------------------------------------
-- binding the routers together
-- connecting router: 0 to router: 2 and vice versa
valid_in_N_2 <= valid_out_S_0;
valid_in_S_0 <= valid_out_N_2;
credit_in_S_0 <= credit_out_N_2;
credit_in_N_2 <= credit_out_S_0;
-------------------
-- connecting router: 1 to router: 3 and vice versa
valid_in_N_3 <= valid_out_S_1;
valid_in_S_1 <= valid_out_N_3;
credit_in_S_1 <= credit_out_N_3;
credit_in_N_3 <= credit_out_S_1;
-------------------

-- connecting router: 0 to router: 1 and vice versa
valid_in_E_0 <= valid_out_W_1;
valid_in_W_1 <= valid_out_E_0;
credit_in_W_1 <= credit_out_E_0;
credit_in_E_0 <= credit_out_W_1;
-------------------
-- connecting router: 2 to router: 3 and vice versa
valid_in_E_2 <= valid_out_W_3;
valid_in_W_3 <= valid_out_E_2;
credit_in_W_3 <= credit_out_E_2;
credit_in_E_2 <= credit_out_W_3;
-------------------
Faulty_S_in0 <= Faulty_N_out2;
Faulty_E_in0 <= Faulty_W_out1;
Faulty_S_in1 <= Faulty_N_out3;
Faulty_W_in1 <= Faulty_E_out0;
Faulty_N_in2 <= Faulty_S_out0;
Faulty_E_in2 <= Faulty_W_out3;
Faulty_N_in3 <= Faulty_S_out1;
Faulty_W_in3 <= Faulty_E_out2;
end;
