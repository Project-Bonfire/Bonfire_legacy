--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated Please do not change!
-- Here are the parameters:
-- 	 network size x:2
-- 	 network size y:2
-- 	 data width:32-- 	 traffic pattern:------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.TB_Package.all;

USE ieee.numeric_std.ALL; 
use IEEE.math_real."ceil";
use IEEE.math_real."log2";

entity tb_network_2x2 is
end tb_network_2x2; 


architecture behavior of tb_network_2x2 is

-- Declaring network component
component network_2x2 is
 generic (DATA_WIDTH: integer := 32; DATA_WIDTH_LV: integer := 11);
port (reset: in  std_logic; 
	clk: in  std_logic; 
	--------------
	RX_L_0: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_0, valid_out_L_0: out std_logic;
	credit_in_L_0, valid_in_L_0: in std_logic;
	TX_L_0: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_1: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_1, valid_out_L_1: out std_logic;
	credit_in_L_1, valid_in_L_1: in std_logic;
	TX_L_1: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_2: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_2, valid_out_L_2: out std_logic;
	credit_in_L_2, valid_in_L_2: in std_logic;
	TX_L_2: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_3: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_3, valid_out_L_3: out std_logic;
	credit_in_L_3, valid_in_L_3: in std_logic;
	TX_L_3: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
    link_faults_0: out std_logic_vector(4 downto 0);
    turn_faults_0: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_0: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_0: in  std_logic_vector(3 downto 0);
    Reconfig_command_0 : in std_logic;

	--------------
    link_faults_1: out std_logic_vector(4 downto 0);
    turn_faults_1: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_1: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_1: in  std_logic_vector(3 downto 0);
    Reconfig_command_1 : in std_logic;

	--------------
    link_faults_2: out std_logic_vector(4 downto 0);
    turn_faults_2: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_2: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_2: in  std_logic_vector(3 downto 0);
    Reconfig_command_2 : in std_logic;

	--------------
    link_faults_3: out std_logic_vector(4 downto 0);
    turn_faults_3: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_3: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_3: in  std_logic_vector(3 downto 0);
    Reconfig_command_3 : in std_logic
            ); 
end component; 
-- Declaring NI component

component NI is
   generic(current_address : integer := 10;   -- the current node's address
           SHMU_address : integer := 0;
           reserved_address : std_logic_vector(29 downto 0) := "000000000000000001111111111111";
           flag_address : std_logic_vector(29 downto 0) :=     "000000000000000010000000000000";  -- reserved address for the memory mapped I/O
           counter_address : std_logic_vector(29 downto 0) :=     "000000000000000010000000000001";
           reconfiguration_address : std_logic_vector(29 downto 0) :=     "000000000000000010000000000010";  -- reserved address for reconfiguration register
           self_diagnosis_address : std_logic_vector(29 downto 0) :=     "000000000000000010000000000011"); -- reserved address for self diagnosis register
   port(clk               : in std_logic;
        reset             : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0);

        -- Flags used by JNIFR and JNIFW instructions
        --NI_read_flag      : out  std_logic;   -- One if the N2P fifo is empty. No read should be performed if one.
        --NI_write_flag      : out  std_logic;  -- One if P2N fifo is full. no write should be performed if one.
        -- interrupt signal: generated evertime a packet is recieved!
        irq_out           : out std_logic;
        -- signals for sending packets to network
        credit_in : in std_logic;
        valid_out: out std_logic;
        TX: out std_logic_vector(31 downto 0);  -- data sent to the NoC
        -- signals for reciving packets from the network
        credit_out : out std_logic;
        valid_in: in std_logic;
        RX: in std_logic_vector(31 downto 0); -- data recieved form the NoC
        -- fault information signals from the router
        link_faults: in std_logic_vector(4 downto 0);
        turn_faults: in std_logic_vector(19 downto 0);

        Rxy_reconf_PE: out  std_logic_vector(7 downto 0);
        Cx_reconf_PE: out  std_logic_vector(3 downto 0);    -- if you are not going to update Cx you should write all ones! (it will be and will the current Cx bits)
        Reconfig_command : out std_logic
  );
end component; --component NI

-- generating bulk signals...
	signal RX_L_0, TX_L_0:  std_logic_vector (31 downto 0);
	signal credit_counter_out_0:  std_logic_vector (1 downto 0);
	signal credit_out_L_0, credit_in_L_0, valid_in_L_0, valid_out_L_0: std_logic;
	signal RX_L_1, TX_L_1:  std_logic_vector (31 downto 0);
	signal credit_counter_out_1:  std_logic_vector (1 downto 0);
	signal credit_out_L_1, credit_in_L_1, valid_in_L_1, valid_out_L_1: std_logic;
	signal RX_L_2, TX_L_2:  std_logic_vector (31 downto 0);
	signal credit_counter_out_2:  std_logic_vector (1 downto 0);
	signal credit_out_L_2, credit_in_L_2, valid_in_L_2, valid_out_L_2: std_logic;
	signal RX_L_3, TX_L_3:  std_logic_vector (31 downto 0);
	signal credit_counter_out_3:  std_logic_vector (1 downto 0);
	signal credit_out_L_3, credit_in_L_3, valid_in_L_3, valid_out_L_3: std_logic;
	signal link_faults_0 : std_logic_vector(4 downto 0);
	signal turn_faults_0 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_0 : std_logic_vector(7 downto 0);
	signal Cx_reconf_PE_0 : std_logic_vector(3 downto 0);
	signal Reconfig_command_0 : std_logic;
	signal link_faults_1 : std_logic_vector(4 downto 0);
	signal turn_faults_1 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_1 : std_logic_vector(7 downto 0);
	signal Cx_reconf_PE_1 : std_logic_vector(3 downto 0);
	signal Reconfig_command_1 : std_logic;
	signal link_faults_2 : std_logic_vector(4 downto 0);
	signal turn_faults_2 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_2 : std_logic_vector(7 downto 0);
	signal Cx_reconf_PE_2 : std_logic_vector(3 downto 0);
	signal Reconfig_command_2 : std_logic;
	signal link_faults_3 : std_logic_vector(4 downto 0);
	signal turn_faults_3 : std_logic_vector(19 downto 0);
	signal Rxy_reconf_PE_3 : std_logic_vector(7 downto 0);
	signal Cx_reconf_PE_3 : std_logic_vector(3 downto 0);
	signal Reconfig_command_3 : std_logic;
	-- NI testing signals
	signal reserved_address :        std_logic_vector(29 downto 0):= "000000000000000001111111111111";
	signal flag_address :            std_logic_vector(29 downto 0):= "000000000000000010000000000000" ; -- reserved address for the memory mapped I/O
	signal counter_address :         std_logic_vector(29 downto 0):= "000000000000000010000000000001";
	signal reconfiguration_address : std_logic_vector(29 downto 0):= "000000000000000010000000000010";  -- reserved address for reconfiguration register
	signal self_diagnosis_address :  std_logic_vector(29 downto 0):= "000000000000000010000000000011";
	signal irq_out_0, irq_out_1, irq_out_2, irq_out_3: std_logic;
	signal test_0, test_1, test_2, test_3: std_logic_vector(31 downto 0);
	signal enable_0, enable_1, enable_2, enable_3: std_logic;
	signal write_byte_enable_0, write_byte_enable_1, write_byte_enable_2, write_byte_enable_3: std_logic_vector(3 downto 0);
	signal address_0, address_1, address_2, address_3: std_logic_vector(31 downto 2);
	signal data_write_0, data_write_1, data_write_2, data_write_3: std_logic_vector(31 downto 0);
	signal data_read_0, data_read_1, data_read_2, data_read_3: std_logic_vector(31 downto 0);
	--------------
	--------------
	constant clk_period : time := 1 ns;
	signal reset, not_reset, clk: std_logic :='0';

begin

   clk_process :process
   begin
        clk <= '0';
        wait for clk_period/2;   
        clk <= '1';
        wait for clk_period/2; 
   end process;

reset <= '1' after 1 ns;
-- instantiating the network
NoC: network_2x2 generic map (DATA_WIDTH  => 32, DATA_WIDTH_LV => 11)
port map (reset, clk, 
	RX_L_0, credit_out_L_0, valid_out_L_0, credit_in_L_0, valid_in_L_0,  TX_L_0, 
	RX_L_1, credit_out_L_1, valid_out_L_1, credit_in_L_1, valid_in_L_1,  TX_L_1, 
	RX_L_2, credit_out_L_2, valid_out_L_2, credit_in_L_2, valid_in_L_2,  TX_L_2, 
	RX_L_3, credit_out_L_3, valid_out_L_3, credit_in_L_3, valid_in_L_3,  TX_L_3, 
	-- should be connected to NI
	link_faults_0, turn_faults_0,	Rxy_reconf_PE_0, Cx_reconf_PE_0, Reconfig_command_0, 
	link_faults_1, turn_faults_1,	Rxy_reconf_PE_1, Cx_reconf_PE_1, Reconfig_command_1, 
	link_faults_2, turn_faults_2,	Rxy_reconf_PE_2, Cx_reconf_PE_2, Reconfig_command_2, 
	link_faults_3, turn_faults_3,	Rxy_reconf_PE_3, Cx_reconf_PE_3, Reconfig_command_3
            ); 
not_reset <= not reset; 

-- connecting the NIs
NI_0: NI 
   generic map(current_address => 0
           ) 
   port map(clk => clk , reset => not_reset , enable => enable_0, 
        write_byte_enable => write_byte_enable_0, 
        address => address_0, 
        data_write => data_write_0, 
        data_read => data_read_0, 
        -- interrupt signal: generated evertime a packet is recieved!
        irq_out => irq_out_0, 
        -- signals for sending packets to network
        credit_in => credit_out_L_0, 
        valid_out => valid_in_L_0,
        TX => RX_L_0, -- data sent to the NoC
        -- signals for reciving packets from the network
        credit_out => credit_in_L_0, 
        valid_in => valid_out_L_0,
        RX => TX_L_0,
        -- fault information signals from the router
        link_faults => link_faults_0, 
        turn_faults => turn_faults_0,

        Rxy_reconf_PE => Rxy_reconf_PE_0, 
        Cx_reconf_PE => Cx_reconf_PE_0,
        Reconfig_command => Reconfig_command_0
  );
NI_1: NI 
   generic map(current_address => 1
           ) 
   port map(clk => clk , reset => not_reset , enable => enable_1, 
        write_byte_enable => write_byte_enable_1, 
        address => address_1, 
        data_write => data_write_1, 
        data_read => data_read_1, 
        -- interrupt signal: generated evertime a packet is recieved!
        irq_out => irq_out_1, 
        -- signals for sending packets to network
        credit_in => credit_out_L_1, 
        valid_out => valid_in_L_1,
        TX => RX_L_1, -- data sent to the NoC
        -- signals for reciving packets from the network
        credit_out => credit_in_L_1, 
        valid_in => valid_out_L_1,
        RX => TX_L_1,
        -- fault information signals from the router
        link_faults => link_faults_1, 
        turn_faults => turn_faults_1,

        Rxy_reconf_PE => Rxy_reconf_PE_1, 
        Cx_reconf_PE => Cx_reconf_PE_1,
        Reconfig_command => Reconfig_command_1
  );
NI_2: NI 
   generic map(current_address => 2
           ) 
   port map(clk => clk , reset => not_reset , enable => enable_2, 
        write_byte_enable => write_byte_enable_2, 
        address => address_2, 
        data_write => data_write_2, 
        data_read => data_read_2, 
        -- interrupt signal: generated evertime a packet is recieved!
        irq_out => irq_out_2, 
        -- signals for sending packets to network
        credit_in => credit_out_L_2, 
        valid_out => valid_in_L_2,
        TX => RX_L_2, -- data sent to the NoC
        -- signals for reciving packets from the network
        credit_out => credit_in_L_2, 
        valid_in => valid_out_L_2,
        RX => TX_L_2,
        -- fault information signals from the router
        link_faults => link_faults_2, 
        turn_faults => turn_faults_2,

        Rxy_reconf_PE => Rxy_reconf_PE_2, 
        Cx_reconf_PE => Cx_reconf_PE_2,
        Reconfig_command => Reconfig_command_2
  );
NI_3: NI 
   generic map(current_address => 3
           ) 
   port map(clk => clk , reset => not_reset , enable => enable_3, 
        write_byte_enable => write_byte_enable_3, 
        address => address_3, 
        data_write => data_write_3, 
        data_read => data_read_3, 
        -- interrupt signal: generated evertime a packet is recieved!
        irq_out => irq_out_3, 
        -- signals for sending packets to network
        credit_in => credit_out_L_3, 
        valid_out => valid_in_L_3,
        TX => RX_L_3, -- data sent to the NoC
        -- signals for reciving packets from the network
        credit_out => credit_in_L_3, 
        valid_in => valid_out_L_3,
        RX => TX_L_3,
        -- fault information signals from the router
        link_faults => link_faults_3, 
        turn_faults => turn_faults_3,

        Rxy_reconf_PE => Rxy_reconf_PE_3, 
        Cx_reconf_PE => Cx_reconf_PE_3,
        Reconfig_command => Reconfig_command_3
  );


-- connecting the packet generators
NI_control(2, 30, 0, 19, 8, 8, 10000 ns, clk,
           -- NI configuration
           reserved_address, flag_address, counter_address, reconfiguration_address, self_diagnosis_address,
           -- NI signals
           enable_0, write_byte_enable_0, address_0, data_write_0, data_read_0, test_0); 

NI_control(2, 30, 1, 20, 8, 8, 10000 ns, clk,
           -- NI configuration
           reserved_address, flag_address, counter_address, reconfiguration_address, self_diagnosis_address,
           -- NI signals
           enable_1, write_byte_enable_1, address_1, data_write_1, data_read_1, test_1); 

NI_control(2, 30, 2, 38, 8, 8, 10000 ns, clk,
           -- NI configuration
           reserved_address, flag_address, counter_address, reconfiguration_address, self_diagnosis_address,
           -- NI signals
           enable_2, write_byte_enable_2, address_2, data_write_2, data_read_2, test_2); 

NI_control(2, 30, 3, 50, 8, 8, 10000 ns, clk,
           -- NI configuration
           reserved_address, flag_address, counter_address, reconfiguration_address, self_diagnosis_address,
           -- NI signals
           enable_3, write_byte_enable_3, address_3, data_write_3, data_read_3, test_3); 



end;
