--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated!
-- Here are the parameters:
-- 	 network size x:4
-- 	 network size y:4
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity network_4x4 is
 generic (DATA_WIDTH: integer := 32);
port (reset: in  std_logic; 
	clk: in  std_logic; 
	--------------
	RX_L_0: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_0, CTS_L_0: out std_logic;
	DRTS_L_0, DCTS_L_0: in std_logic;
	TX_L_0: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_1: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_1, CTS_L_1: out std_logic;
	DRTS_L_1, DCTS_L_1: in std_logic;
	TX_L_1: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_2: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_2, CTS_L_2: out std_logic;
	DRTS_L_2, DCTS_L_2: in std_logic;
	TX_L_2: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_3: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_3, CTS_L_3: out std_logic;
	DRTS_L_3, DCTS_L_3: in std_logic;
	TX_L_3: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_4: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_4, CTS_L_4: out std_logic;
	DRTS_L_4, DCTS_L_4: in std_logic;
	TX_L_4: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_5: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_5, CTS_L_5: out std_logic;
	DRTS_L_5, DCTS_L_5: in std_logic;
	TX_L_5: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_6: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_6, CTS_L_6: out std_logic;
	DRTS_L_6, DCTS_L_6: in std_logic;
	TX_L_6: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_7: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_7, CTS_L_7: out std_logic;
	DRTS_L_7, DCTS_L_7: in std_logic;
	TX_L_7: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_8: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_8, CTS_L_8: out std_logic;
	DRTS_L_8, DCTS_L_8: in std_logic;
	TX_L_8: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_9: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_9, CTS_L_9: out std_logic;
	DRTS_L_9, DCTS_L_9: in std_logic;
	TX_L_9: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_10: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_10, CTS_L_10: out std_logic;
	DRTS_L_10, DCTS_L_10: in std_logic;
	TX_L_10: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_11: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_11, CTS_L_11: out std_logic;
	DRTS_L_11, DCTS_L_11: in std_logic;
	TX_L_11: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_12: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_12, CTS_L_12: out std_logic;
	DRTS_L_12, DCTS_L_12: in std_logic;
	TX_L_12: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_13: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_13, CTS_L_13: out std_logic;
	DRTS_L_13, DCTS_L_13: in std_logic;
	TX_L_13: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_14: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_14, CTS_L_14: out std_logic;
	DRTS_L_14, DCTS_L_14: in std_logic;
	TX_L_14: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_15: in std_logic_vector (DATA_WIDTH-1 downto 0);
	RTS_L_15, CTS_L_15: out std_logic;
	DRTS_L_15, DCTS_L_15: in std_logic;
	TX_L_15: out std_logic_vector (DATA_WIDTH-1 downto 0)
            ); 
end network_4x4; 


architecture behavior of network_4x4 is

-- Declaring router component
component router is
 generic (
        DATA_WIDTH: integer := 32;
        current_address : integer := 5;
        Rxy_rst : integer := 60;
        Cx_rst : integer := 15
    );
    port (
    reset, clk: in std_logic;
    DCTS_N, DCTS_E, DCTS_w, DCTS_S, DCTS_L: in std_logic;
    DRTS_N, DRTS_E, DRTS_W, DRTS_S, DRTS_L: in std_logic;
    RX_N, RX_E, RX_W, RX_S, RX_L : in std_logic_vector (DATA_WIDTH-1 downto 0);
    RTS_N, RTS_E, RTS_W, RTS_S, RTS_L: out std_logic;
    CTS_N, CTS_E, CTS_w, CTS_S, CTS_L: out std_logic;
    TX_N, TX_E, TX_W, TX_S, TX_L: out std_logic_vector (DATA_WIDTH-1 downto 0));
end component; 

-- generating bulk signals. not all of them are used in the design...
	signal DCTS_N_0, DCTS_E_0, DCTS_w_0, DCTS_S_0: std_logic;
	signal DCTS_N_1, DCTS_E_1, DCTS_w_1, DCTS_S_1: std_logic;
	signal DCTS_N_2, DCTS_E_2, DCTS_w_2, DCTS_S_2: std_logic;
	signal DCTS_N_3, DCTS_E_3, DCTS_w_3, DCTS_S_3: std_logic;
	signal DCTS_N_4, DCTS_E_4, DCTS_w_4, DCTS_S_4: std_logic;
	signal DCTS_N_5, DCTS_E_5, DCTS_w_5, DCTS_S_5: std_logic;
	signal DCTS_N_6, DCTS_E_6, DCTS_w_6, DCTS_S_6: std_logic;
	signal DCTS_N_7, DCTS_E_7, DCTS_w_7, DCTS_S_7: std_logic;
	signal DCTS_N_8, DCTS_E_8, DCTS_w_8, DCTS_S_8: std_logic;
	signal DCTS_N_9, DCTS_E_9, DCTS_w_9, DCTS_S_9: std_logic;
	signal DCTS_N_10, DCTS_E_10, DCTS_w_10, DCTS_S_10: std_logic;
	signal DCTS_N_11, DCTS_E_11, DCTS_w_11, DCTS_S_11: std_logic;
	signal DCTS_N_12, DCTS_E_12, DCTS_w_12, DCTS_S_12: std_logic;
	signal DCTS_N_13, DCTS_E_13, DCTS_w_13, DCTS_S_13: std_logic;
	signal DCTS_N_14, DCTS_E_14, DCTS_w_14, DCTS_S_14: std_logic;
	signal DCTS_N_15, DCTS_E_15, DCTS_w_15, DCTS_S_15: std_logic;

	signal DRTS_N_0, DRTS_E_0, DRTS_W_0, DRTS_S_0: std_logic;
	signal DRTS_N_1, DRTS_E_1, DRTS_W_1, DRTS_S_1: std_logic;
	signal DRTS_N_2, DRTS_E_2, DRTS_W_2, DRTS_S_2: std_logic;
	signal DRTS_N_3, DRTS_E_3, DRTS_W_3, DRTS_S_3: std_logic;
	signal DRTS_N_4, DRTS_E_4, DRTS_W_4, DRTS_S_4: std_logic;
	signal DRTS_N_5, DRTS_E_5, DRTS_W_5, DRTS_S_5: std_logic;
	signal DRTS_N_6, DRTS_E_6, DRTS_W_6, DRTS_S_6: std_logic;
	signal DRTS_N_7, DRTS_E_7, DRTS_W_7, DRTS_S_7: std_logic;
	signal DRTS_N_8, DRTS_E_8, DRTS_W_8, DRTS_S_8: std_logic;
	signal DRTS_N_9, DRTS_E_9, DRTS_W_9, DRTS_S_9: std_logic;
	signal DRTS_N_10, DRTS_E_10, DRTS_W_10, DRTS_S_10: std_logic;
	signal DRTS_N_11, DRTS_E_11, DRTS_W_11, DRTS_S_11: std_logic;
	signal DRTS_N_12, DRTS_E_12, DRTS_W_12, DRTS_S_12: std_logic;
	signal DRTS_N_13, DRTS_E_13, DRTS_W_13, DRTS_S_13: std_logic;
	signal DRTS_N_14, DRTS_E_14, DRTS_W_14, DRTS_S_14: std_logic;
	signal DRTS_N_15, DRTS_E_15, DRTS_W_15, DRTS_S_15: std_logic;

	signal RX_N_0, RX_E_0, RX_W_0, RX_S_0 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_1, RX_E_1, RX_W_1, RX_S_1 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_2, RX_E_2, RX_W_2, RX_S_2 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_3, RX_E_3, RX_W_3, RX_S_3 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_4, RX_E_4, RX_W_4, RX_S_4 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_5, RX_E_5, RX_W_5, RX_S_5 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_6, RX_E_6, RX_W_6, RX_S_6 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_7, RX_E_7, RX_W_7, RX_S_7 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_8, RX_E_8, RX_W_8, RX_S_8 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_9, RX_E_9, RX_W_9, RX_S_9 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_10, RX_E_10, RX_W_10, RX_S_10 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_11, RX_E_11, RX_W_11, RX_S_11 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_12, RX_E_12, RX_W_12, RX_S_12 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_13, RX_E_13, RX_W_13, RX_S_13 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_14, RX_E_14, RX_W_14, RX_S_14 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_15, RX_E_15, RX_W_15, RX_S_15 : std_logic_vector (DATA_WIDTH-1 downto 0);

	signal CTS_N_0, CTS_E_0, CTS_w_0, CTS_S_0: std_logic;
	signal CTS_N_1, CTS_E_1, CTS_w_1, CTS_S_1: std_logic;
	signal CTS_N_2, CTS_E_2, CTS_w_2, CTS_S_2: std_logic;
	signal CTS_N_3, CTS_E_3, CTS_w_3, CTS_S_3: std_logic;
	signal CTS_N_4, CTS_E_4, CTS_w_4, CTS_S_4: std_logic;
	signal CTS_N_5, CTS_E_5, CTS_w_5, CTS_S_5: std_logic;
	signal CTS_N_6, CTS_E_6, CTS_w_6, CTS_S_6: std_logic;
	signal CTS_N_7, CTS_E_7, CTS_w_7, CTS_S_7: std_logic;
	signal CTS_N_8, CTS_E_8, CTS_w_8, CTS_S_8: std_logic;
	signal CTS_N_9, CTS_E_9, CTS_w_9, CTS_S_9: std_logic;
	signal CTS_N_10, CTS_E_10, CTS_w_10, CTS_S_10: std_logic;
	signal CTS_N_11, CTS_E_11, CTS_w_11, CTS_S_11: std_logic;
	signal CTS_N_12, CTS_E_12, CTS_w_12, CTS_S_12: std_logic;
	signal CTS_N_13, CTS_E_13, CTS_w_13, CTS_S_13: std_logic;
	signal CTS_N_14, CTS_E_14, CTS_w_14, CTS_S_14: std_logic;
	signal CTS_N_15, CTS_E_15, CTS_w_15, CTS_S_15: std_logic;

	signal RTS_N_0, RTS_E_0, RTS_W_0, RTS_S_0: std_logic;
	signal RTS_N_1, RTS_E_1, RTS_W_1, RTS_S_1: std_logic;
	signal RTS_N_2, RTS_E_2, RTS_W_2, RTS_S_2: std_logic;
	signal RTS_N_3, RTS_E_3, RTS_W_3, RTS_S_3: std_logic;
	signal RTS_N_4, RTS_E_4, RTS_W_4, RTS_S_4: std_logic;
	signal RTS_N_5, RTS_E_5, RTS_W_5, RTS_S_5: std_logic;
	signal RTS_N_6, RTS_E_6, RTS_W_6, RTS_S_6: std_logic;
	signal RTS_N_7, RTS_E_7, RTS_W_7, RTS_S_7: std_logic;
	signal RTS_N_8, RTS_E_8, RTS_W_8, RTS_S_8: std_logic;
	signal RTS_N_9, RTS_E_9, RTS_W_9, RTS_S_9: std_logic;
	signal RTS_N_10, RTS_E_10, RTS_W_10, RTS_S_10: std_logic;
	signal RTS_N_11, RTS_E_11, RTS_W_11, RTS_S_11: std_logic;
	signal RTS_N_12, RTS_E_12, RTS_W_12, RTS_S_12: std_logic;
	signal RTS_N_13, RTS_E_13, RTS_W_13, RTS_S_13: std_logic;
	signal RTS_N_14, RTS_E_14, RTS_W_14, RTS_S_14: std_logic;
	signal RTS_N_15, RTS_E_15, RTS_W_15, RTS_S_15: std_logic;

	signal TX_N_0, TX_E_0, TX_W_0, TX_S_0 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_1, TX_E_1, TX_W_1, TX_S_1 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_2, TX_E_2, TX_W_2, TX_S_2 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_3, TX_E_3, TX_W_3, TX_S_3 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_4, TX_E_4, TX_W_4, TX_S_4 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_5, TX_E_5, TX_W_5, TX_S_5 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_6, TX_E_6, TX_W_6, TX_S_6 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_7, TX_E_7, TX_W_7, TX_S_7 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_8, TX_E_8, TX_W_8, TX_S_8 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_9, TX_E_9, TX_W_9, TX_S_9 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_10, TX_E_10, TX_W_10, TX_S_10 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_11, TX_E_11, TX_W_11, TX_S_11 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_12, TX_E_12, TX_W_12, TX_S_12 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_13, TX_E_13, TX_W_13, TX_S_13 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_14, TX_E_14, TX_W_14, TX_S_14 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_15, TX_E_15, TX_W_15, TX_S_15 : std_logic_vector (DATA_WIDTH-1 downto 0);
begin

-- instantiating the routers
R_0: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>0, Rxy_rst => 60, Cx_rst => 10)
PORT MAP (reset, clk, 
	DCTS_N_0, DCTS_E_0, DCTS_W_0, DCTS_S_0, DCTS_L_0,
	DRTS_N_0, DRTS_E_0, DRTS_W_0, DRTS_S_0, DRTS_L_0,
	RX_N_0, RX_E_0, RX_W_0, RX_S_0, RX_L_0,
	RTS_N_0, RTS_E_0, RTS_W_0, RTS_S_0, RTS_L_0,
	CTS_N_0, CTS_E_0, CTS_w_0, CTS_S_0, CTS_L_0,
	TX_N_0, TX_E_0, TX_W_0, TX_S_0, TX_L_0); 

R_1: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>1, Rxy_rst => 60, Cx_rst => 14)
PORT MAP (reset, clk, 
	DCTS_N_1, DCTS_E_1, DCTS_W_1, DCTS_S_1, DCTS_L_1,
	DRTS_N_1, DRTS_E_1, DRTS_W_1, DRTS_S_1, DRTS_L_1,
	RX_N_1, RX_E_1, RX_W_1, RX_S_1, RX_L_1,
	RTS_N_1, RTS_E_1, RTS_W_1, RTS_S_1, RTS_L_1,
	CTS_N_1, CTS_E_1, CTS_w_1, CTS_S_1, CTS_L_1,
	TX_N_1, TX_E_1, TX_W_1, TX_S_1, TX_L_1); 

R_2: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>2, Rxy_rst => 60, Cx_rst => 14)
PORT MAP (reset, clk, 
	DCTS_N_2, DCTS_E_2, DCTS_W_2, DCTS_S_2, DCTS_L_2,
	DRTS_N_2, DRTS_E_2, DRTS_W_2, DRTS_S_2, DRTS_L_2,
	RX_N_2, RX_E_2, RX_W_2, RX_S_2, RX_L_2,
	RTS_N_2, RTS_E_2, RTS_W_2, RTS_S_2, RTS_L_2,
	CTS_N_2, CTS_E_2, CTS_w_2, CTS_S_2, CTS_L_2,
	TX_N_2, TX_E_2, TX_W_2, TX_S_2, TX_L_2); 

R_3: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>3, Rxy_rst => 60, Cx_rst => 12)
PORT MAP (reset, clk, 
	DCTS_N_3, DCTS_E_3, DCTS_W_3, DCTS_S_3, DCTS_L_3,
	DRTS_N_3, DRTS_E_3, DRTS_W_3, DRTS_S_3, DRTS_L_3,
	RX_N_3, RX_E_3, RX_W_3, RX_S_3, RX_L_3,
	RTS_N_3, RTS_E_3, RTS_W_3, RTS_S_3, RTS_L_3,
	CTS_N_3, CTS_E_3, CTS_w_3, CTS_S_3, CTS_L_3,
	TX_N_3, TX_E_3, TX_W_3, TX_S_3, TX_L_3); 

R_4: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>4, Rxy_rst => 60, Cx_rst => 11)
PORT MAP (reset, clk, 
	DCTS_N_4, DCTS_E_4, DCTS_W_4, DCTS_S_4, DCTS_L_4,
	DRTS_N_4, DRTS_E_4, DRTS_W_4, DRTS_S_4, DRTS_L_4,
	RX_N_4, RX_E_4, RX_W_4, RX_S_4, RX_L_4,
	RTS_N_4, RTS_E_4, RTS_W_4, RTS_S_4, RTS_L_4,
	CTS_N_4, CTS_E_4, CTS_w_4, CTS_S_4, CTS_L_4,
	TX_N_4, TX_E_4, TX_W_4, TX_S_4, TX_L_4); 

R_5: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>5, Rxy_rst => 60, Cx_rst => 15)
PORT MAP (reset, clk, 
	DCTS_N_5, DCTS_E_5, DCTS_W_5, DCTS_S_5, DCTS_L_5,
	DRTS_N_5, DRTS_E_5, DRTS_W_5, DRTS_S_5, DRTS_L_5,
	RX_N_5, RX_E_5, RX_W_5, RX_S_5, RX_L_5,
	RTS_N_5, RTS_E_5, RTS_W_5, RTS_S_5, RTS_L_5,
	CTS_N_5, CTS_E_5, CTS_w_5, CTS_S_5, CTS_L_5,
	TX_N_5, TX_E_5, TX_W_5, TX_S_5, TX_L_5); 

R_6: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>6, Rxy_rst => 60, Cx_rst => 15)
PORT MAP (reset, clk, 
	DCTS_N_6, DCTS_E_6, DCTS_W_6, DCTS_S_6, DCTS_L_6,
	DRTS_N_6, DRTS_E_6, DRTS_W_6, DRTS_S_6, DRTS_L_6,
	RX_N_6, RX_E_6, RX_W_6, RX_S_6, RX_L_6,
	RTS_N_6, RTS_E_6, RTS_W_6, RTS_S_6, RTS_L_6,
	CTS_N_6, CTS_E_6, CTS_w_6, CTS_S_6, CTS_L_6,
	TX_N_6, TX_E_6, TX_W_6, TX_S_6, TX_L_6); 

R_7: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>7, Rxy_rst => 60, Cx_rst => 13)
PORT MAP (reset, clk, 
	DCTS_N_7, DCTS_E_7, DCTS_W_7, DCTS_S_7, DCTS_L_7,
	DRTS_N_7, DRTS_E_7, DRTS_W_7, DRTS_S_7, DRTS_L_7,
	RX_N_7, RX_E_7, RX_W_7, RX_S_7, RX_L_7,
	RTS_N_7, RTS_E_7, RTS_W_7, RTS_S_7, RTS_L_7,
	CTS_N_7, CTS_E_7, CTS_w_7, CTS_S_7, CTS_L_7,
	TX_N_7, TX_E_7, TX_W_7, TX_S_7, TX_L_7); 

R_8: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>8, Rxy_rst => 60, Cx_rst => 11)
PORT MAP (reset, clk, 
	DCTS_N_8, DCTS_E_8, DCTS_W_8, DCTS_S_8, DCTS_L_8,
	DRTS_N_8, DRTS_E_8, DRTS_W_8, DRTS_S_8, DRTS_L_8,
	RX_N_8, RX_E_8, RX_W_8, RX_S_8, RX_L_8,
	RTS_N_8, RTS_E_8, RTS_W_8, RTS_S_8, RTS_L_8,
	CTS_N_8, CTS_E_8, CTS_w_8, CTS_S_8, CTS_L_8,
	TX_N_8, TX_E_8, TX_W_8, TX_S_8, TX_L_8); 

R_9: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>9, Rxy_rst => 60, Cx_rst => 15)
PORT MAP (reset, clk, 
	DCTS_N_9, DCTS_E_9, DCTS_W_9, DCTS_S_9, DCTS_L_9,
	DRTS_N_9, DRTS_E_9, DRTS_W_9, DRTS_S_9, DRTS_L_9,
	RX_N_9, RX_E_9, RX_W_9, RX_S_9, RX_L_9,
	RTS_N_9, RTS_E_9, RTS_W_9, RTS_S_9, RTS_L_9,
	CTS_N_9, CTS_E_9, CTS_w_9, CTS_S_9, CTS_L_9,
	TX_N_9, TX_E_9, TX_W_9, TX_S_9, TX_L_9); 

R_10: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>10, Rxy_rst => 60, Cx_rst => 15)
PORT MAP (reset, clk, 
	DCTS_N_10, DCTS_E_10, DCTS_W_10, DCTS_S_10, DCTS_L_10,
	DRTS_N_10, DRTS_E_10, DRTS_W_10, DRTS_S_10, DRTS_L_10,
	RX_N_10, RX_E_10, RX_W_10, RX_S_10, RX_L_10,
	RTS_N_10, RTS_E_10, RTS_W_10, RTS_S_10, RTS_L_10,
	CTS_N_10, CTS_E_10, CTS_w_10, CTS_S_10, CTS_L_10,
	TX_N_10, TX_E_10, TX_W_10, TX_S_10, TX_L_10); 

R_11: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>11, Rxy_rst => 60, Cx_rst => 13)
PORT MAP (reset, clk, 
	DCTS_N_11, DCTS_E_11, DCTS_W_11, DCTS_S_11, DCTS_L_11,
	DRTS_N_11, DRTS_E_11, DRTS_W_11, DRTS_S_11, DRTS_L_11,
	RX_N_11, RX_E_11, RX_W_11, RX_S_11, RX_L_11,
	RTS_N_11, RTS_E_11, RTS_W_11, RTS_S_11, RTS_L_11,
	CTS_N_11, CTS_E_11, CTS_w_11, CTS_S_11, CTS_L_11,
	TX_N_11, TX_E_11, TX_W_11, TX_S_11, TX_L_11); 

R_12: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>12, Rxy_rst => 60, Cx_rst => 3)
PORT MAP (reset, clk, 
	DCTS_N_12, DCTS_E_12, DCTS_W_12, DCTS_S_12, DCTS_L_12,
	DRTS_N_12, DRTS_E_12, DRTS_W_12, DRTS_S_12, DRTS_L_12,
	RX_N_12, RX_E_12, RX_W_12, RX_S_12, RX_L_12,
	RTS_N_12, RTS_E_12, RTS_W_12, RTS_S_12, RTS_L_12,
	CTS_N_12, CTS_E_12, CTS_w_12, CTS_S_12, CTS_L_12,
	TX_N_12, TX_E_12, TX_W_12, TX_S_12, TX_L_12); 

R_13: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>13, Rxy_rst => 60, Cx_rst => 7)
PORT MAP (reset, clk, 
	DCTS_N_13, DCTS_E_13, DCTS_W_13, DCTS_S_13, DCTS_L_13,
	DRTS_N_13, DRTS_E_13, DRTS_W_13, DRTS_S_13, DRTS_L_13,
	RX_N_13, RX_E_13, RX_W_13, RX_S_13, RX_L_13,
	RTS_N_13, RTS_E_13, RTS_W_13, RTS_S_13, RTS_L_13,
	CTS_N_13, CTS_E_13, CTS_w_13, CTS_S_13, CTS_L_13,
	TX_N_13, TX_E_13, TX_W_13, TX_S_13, TX_L_13); 

R_14: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>14, Rxy_rst => 60, Cx_rst => 7)
PORT MAP (reset, clk, 
	DCTS_N_14, DCTS_E_14, DCTS_W_14, DCTS_S_14, DCTS_L_14,
	DRTS_N_14, DRTS_E_14, DRTS_W_14, DRTS_S_14, DRTS_L_14,
	RX_N_14, RX_E_14, RX_W_14, RX_S_14, RX_L_14,
	RTS_N_14, RTS_E_14, RTS_W_14, RTS_S_14, RTS_L_14,
	CTS_N_14, CTS_E_14, CTS_w_14, CTS_S_14, CTS_L_14,
	TX_N_14, TX_E_14, TX_W_14, TX_S_14, TX_L_14); 

R_15: router generic map (DATA_WIDTH  => DATA_WIDTH, current_address=>15, Rxy_rst => 60, Cx_rst => 5)
PORT MAP (reset, clk, 
	DCTS_N_15, DCTS_E_15, DCTS_W_15, DCTS_S_15, DCTS_L_15,
	DRTS_N_15, DRTS_E_15, DRTS_W_15, DRTS_S_15, DRTS_L_15,
	RX_N_15, RX_E_15, RX_W_15, RX_S_15, RX_L_15,
	RTS_N_15, RTS_E_15, RTS_W_15, RTS_S_15, RTS_L_15,
	CTS_N_15, CTS_E_15, CTS_w_15, CTS_S_15, CTS_L_15,
	TX_N_15, TX_E_15, TX_W_15, TX_S_15, TX_L_15); 

-- binding the routers together
-- vertical ins/outs
-- connecting router: 0 to router: 4 and vice versa
RX_N_4<= TX_S_0;
RX_S_0<= TX_N_4;
DRTS_N_4 <= RTS_S_0;
DCTS_S_0 <= CTS_N_4;
DRTS_S_0 <= RTS_N_4;
DCTS_N_4 <= CTS_S_0;
-------------------
-- connecting router: 1 to router: 5 and vice versa
RX_N_5<= TX_S_1;
RX_S_1<= TX_N_5;
DRTS_N_5 <= RTS_S_1;
DCTS_S_1 <= CTS_N_5;
DRTS_S_1 <= RTS_N_5;
DCTS_N_5 <= CTS_S_1;
-------------------
-- connecting router: 2 to router: 6 and vice versa
RX_N_6<= TX_S_2;
RX_S_2<= TX_N_6;
DRTS_N_6 <= RTS_S_2;
DCTS_S_2 <= CTS_N_6;
DRTS_S_2 <= RTS_N_6;
DCTS_N_6 <= CTS_S_2;
-------------------
-- connecting router: 3 to router: 7 and vice versa
RX_N_7<= TX_S_3;
RX_S_3<= TX_N_7;
DRTS_N_7 <= RTS_S_3;
DCTS_S_3 <= CTS_N_7;
DRTS_S_3 <= RTS_N_7;
DCTS_N_7 <= CTS_S_3;
-------------------
-- connecting router: 4 to router: 8 and vice versa
RX_N_8<= TX_S_4;
RX_S_4<= TX_N_8;
DRTS_N_8 <= RTS_S_4;
DCTS_S_4 <= CTS_N_8;
DRTS_S_4 <= RTS_N_8;
DCTS_N_8 <= CTS_S_4;
-------------------
-- connecting router: 5 to router: 9 and vice versa
RX_N_9<= TX_S_5;
RX_S_5<= TX_N_9;
DRTS_N_9 <= RTS_S_5;
DCTS_S_5 <= CTS_N_9;
DRTS_S_5 <= RTS_N_9;
DCTS_N_9 <= CTS_S_5;
-------------------
-- connecting router: 6 to router: 10 and vice versa
RX_N_10<= TX_S_6;
RX_S_6<= TX_N_10;
DRTS_N_10 <= RTS_S_6;
DCTS_S_6 <= CTS_N_10;
DRTS_S_6 <= RTS_N_10;
DCTS_N_10 <= CTS_S_6;
-------------------
-- connecting router: 7 to router: 11 and vice versa
RX_N_11<= TX_S_7;
RX_S_7<= TX_N_11;
DRTS_N_11 <= RTS_S_7;
DCTS_S_7 <= CTS_N_11;
DRTS_S_7 <= RTS_N_11;
DCTS_N_11 <= CTS_S_7;
-------------------
-- connecting router: 8 to router: 12 and vice versa
RX_N_12<= TX_S_8;
RX_S_8<= TX_N_12;
DRTS_N_12 <= RTS_S_8;
DCTS_S_8 <= CTS_N_12;
DRTS_S_8 <= RTS_N_12;
DCTS_N_12 <= CTS_S_8;
-------------------
-- connecting router: 9 to router: 13 and vice versa
RX_N_13<= TX_S_9;
RX_S_9<= TX_N_13;
DRTS_N_13 <= RTS_S_9;
DCTS_S_9 <= CTS_N_13;
DRTS_S_9 <= RTS_N_13;
DCTS_N_13 <= CTS_S_9;
-------------------
-- connecting router: 10 to router: 14 and vice versa
RX_N_14<= TX_S_10;
RX_S_10<= TX_N_14;
DRTS_N_14 <= RTS_S_10;
DCTS_S_10 <= CTS_N_14;
DRTS_S_10 <= RTS_N_14;
DCTS_N_14 <= CTS_S_10;
-------------------
-- connecting router: 11 to router: 15 and vice versa
RX_N_15<= TX_S_11;
RX_S_11<= TX_N_15;
DRTS_N_15 <= RTS_S_11;
DCTS_S_11 <= CTS_N_15;
DRTS_S_11 <= RTS_N_15;
DCTS_N_15 <= CTS_S_11;
-------------------

-- horizontal ins/outs
-- connecting router: 0 to router: 1 and vice versa
RX_E_0 <= TX_W_1;
RX_W_1 <= TX_E_0;
DRTS_E_0 <= RTS_W_1;
DCTS_W_1 <= CTS_E_0;
DRTS_W_1 <= RTS_E_0;
DCTS_E_0 <= CTS_W_1;
-------------------
-- connecting router: 1 to router: 2 and vice versa
RX_E_1 <= TX_W_2;
RX_W_2 <= TX_E_1;
DRTS_E_1 <= RTS_W_2;
DCTS_W_2 <= CTS_E_1;
DRTS_W_2 <= RTS_E_1;
DCTS_E_1 <= CTS_W_2;
-------------------
-- connecting router: 2 to router: 3 and vice versa
RX_E_2 <= TX_W_3;
RX_W_3 <= TX_E_2;
DRTS_E_2 <= RTS_W_3;
DCTS_W_3 <= CTS_E_2;
DRTS_W_3 <= RTS_E_2;
DCTS_E_2 <= CTS_W_3;
-------------------
-- connecting router: 4 to router: 5 and vice versa
RX_E_4 <= TX_W_5;
RX_W_5 <= TX_E_4;
DRTS_E_4 <= RTS_W_5;
DCTS_W_5 <= CTS_E_4;
DRTS_W_5 <= RTS_E_4;
DCTS_E_4 <= CTS_W_5;
-------------------
-- connecting router: 5 to router: 6 and vice versa
RX_E_5 <= TX_W_6;
RX_W_6 <= TX_E_5;
DRTS_E_5 <= RTS_W_6;
DCTS_W_6 <= CTS_E_5;
DRTS_W_6 <= RTS_E_5;
DCTS_E_5 <= CTS_W_6;
-------------------
-- connecting router: 6 to router: 7 and vice versa
RX_E_6 <= TX_W_7;
RX_W_7 <= TX_E_6;
DRTS_E_6 <= RTS_W_7;
DCTS_W_7 <= CTS_E_6;
DRTS_W_7 <= RTS_E_6;
DCTS_E_6 <= CTS_W_7;
-------------------
-- connecting router: 8 to router: 9 and vice versa
RX_E_8 <= TX_W_9;
RX_W_9 <= TX_E_8;
DRTS_E_8 <= RTS_W_9;
DCTS_W_9 <= CTS_E_8;
DRTS_W_9 <= RTS_E_8;
DCTS_E_8 <= CTS_W_9;
-------------------
-- connecting router: 9 to router: 10 and vice versa
RX_E_9 <= TX_W_10;
RX_W_10 <= TX_E_9;
DRTS_E_9 <= RTS_W_10;
DCTS_W_10 <= CTS_E_9;
DRTS_W_10 <= RTS_E_9;
DCTS_E_9 <= CTS_W_10;
-------------------
-- connecting router: 10 to router: 11 and vice versa
RX_E_10 <= TX_W_11;
RX_W_11 <= TX_E_10;
DRTS_E_10 <= RTS_W_11;
DCTS_W_11 <= CTS_E_10;
DRTS_W_11 <= RTS_E_10;
DCTS_E_10 <= CTS_W_11;
-------------------
-- connecting router: 12 to router: 13 and vice versa
RX_E_12 <= TX_W_13;
RX_W_13 <= TX_E_12;
DRTS_E_12 <= RTS_W_13;
DCTS_W_13 <= CTS_E_12;
DRTS_W_13 <= RTS_E_12;
DCTS_E_12 <= CTS_W_13;
-------------------
-- connecting router: 13 to router: 14 and vice versa
RX_E_13 <= TX_W_14;
RX_W_14 <= TX_E_13;
DRTS_E_13 <= RTS_W_14;
DCTS_W_14 <= CTS_E_13;
DRTS_W_14 <= RTS_E_13;
DCTS_E_13 <= CTS_W_14;
-------------------
-- connecting router: 14 to router: 15 and vice versa
RX_E_14 <= TX_W_15;
RX_W_15 <= TX_E_14;
DRTS_E_14 <= RTS_W_15;
DCTS_W_15 <= CTS_E_14;
DRTS_W_15 <= RTS_E_14;
DCTS_E_14 <= CTS_W_15;
-------------------
end;

