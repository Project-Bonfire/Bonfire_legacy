--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated!
-- Here are the parameters:
-- 	 network size x: 2
-- 	 network size y: 2
-- 	 Data width: 32
-- 	 Parity: False
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.numeric_std.ALL;
use work.component_pack.all;

entity toppest_module is
 generic (DATA_WIDTH: integer := 32;
          -- DATA_WIDTH_LV: integer := 11;
          memory_type : string :=
--             "TRI_PORT_X"
           --   "DUAL_PORT_"
           --   "ALTERA_LPM"
               "XILINX_16X"
      );

port (
      reset: in  std_logic;
      clk: in  std_logic;

      -- IJTAG network for fault injection and checker status monitoring
      TCK         : in std_logic;
      RST         : in std_logic;
      SEL         : in std_logic;
      SI          : in std_logic;
      SE          : in std_logic;
      UE          : in std_logic;
      CE          : in std_logic;
      SO          : out std_logic;
      toF         : out std_logic;
      toC         : out std_logic;

      -- GPIO for Node 0
      GPIO_out: out  std_logic_vector(15 downto 0);
      GPIO_in: in  std_logic_vector(14 downto 0);
--      GPIO_in: in  std_logic_vector(21 downto 15); --not enough inputs

      -- UART for all Plasmas
      uart_write_0  : out std_logic;
      uart_read_0   : in std_logic;
      uart_write_1  : out std_logic;
      uart_read_1   : in std_logic;
      uart_write_2  : out std_logic;
      uart_read_2   : in std_logic;
      uart_write_3  : out std_logic;
      uart_read_3   : in std_logic
    );

end toppest_module;



architecture behavior of toppest_module is
signal clk1_noc, clk2_ijtag : std_logic;

begin


       noc2x2_inst: entity work.network_2x2_with_PE
       generic map (
        DATA_WIDTH => DATA_WIDTH,
        DATA_WIDTH_LV => 0, --UNUSED
        memory_type => memory_type
       )
       port map (
        reset => reset,
        clk => clk1_noc,

        TCK => clk2_ijtag,
        RST => RST,
        SEL => SEL,
        SI => SI,
        SE => SE,
        UE => UE,
        CE => CE,
        SO => SO,
        toF => toF,
        toC => toC,

        GPIO_out => GPIO_out,
        GPIO_in => "0000000" & GPIO_in, --switch(0) == GPIO_in(0) ...


        uart_write_0 => uart_write_0,
        uart_read_0 => uart_read_0,
        uart_write_1 => uart_write_1,
        uart_read_1 => uart_read_1,
        uart_write_2 => uart_write_2,
        uart_read_2 => uart_read_2,
        uart_write_3 => uart_write_3,
        uart_read_3 => uart_read_3
          );



       clk_gen: entity work.clk_wiz_0
       port map (
          --in:
          clk_in1       => clk,

          --out:
          clk1_noc       => clk1_noc,
          clk2_ijtag     => clk2_ijtag);

end;
