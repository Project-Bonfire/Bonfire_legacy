--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated Please do not change!
-- Here are the parameters:
-- 	 network size x:2
-- 	 network size y:2
-- 	 data width:32-- 	 traffic pattern:------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--use work.TB_Package.all;
use work.mlite_pack.all;

USE ieee.numeric_std.ALL;
--use IEEE.math_real."ceil";
--use IEEE.math_real."log2";

entity tb_network_2x2 is
end tb_network_2x2;


architecture behavior of tb_network_2x2 is

constant fcXS : std_logic_vector(0 to 3) := "1011";
constant fcXN : std_logic_vector(0 to 3) := "1010";
constant RAMDataSize : positive := 32;
constant RAMAddrSize : positive := 12;
constant path : string(1 to 12) := "Testbenches/"; --uncomment this if you are SIMULATING in MODELSIM, or if you're synthesizing.
-- constant path : string(positive range <>) := "/home/tsotne/ownCloud/git/Bonfire_sim/Bonfire/RTL/Chip_Designs/IMMORTAL_Chip_2017/Testbenches/"; --used only for Vivado similation. Tsotnes PC.

-- Declaring network component
component network_2x2_with_PE is
 generic (DATA_WIDTH: integer := 32; DATA_WIDTH_LV: integer := 11);
port (reset: in  std_logic;
      clk: in  std_logic;

      -- IJTAG network for fault injection and checker status monitoring
      TCK         : in std_logic;
      RST         : in std_logic;
      SEL         : in std_logic;
      SI          : in std_logic;
      SE          : in std_logic;
      UE          : in std_logic;
      CE          : in std_logic;
      SO          : out std_logic;
      toF         : out std_logic;
      toC         : out std_logic;

      -- GPIO for Node 0
      GPIO_out: out  std_logic_vector(15 downto 0);
      GPIO_in: in  std_logic_vector(21 downto 0);
           -- UART for all Plasmas
      uart_write_0  : out std_logic;
      uart_read_0   : in std_logic;
      uart_write_1  : out std_logic;
      uart_read_1   : in std_logic;
      uart_write_2  : out std_logic;
      uart_read_2   : in std_logic;
      uart_write_3  : out std_logic;
      uart_read_3   : in std_logic;

      -- Monitor connections
      temperature_control   : out std_logic_vector(2 downto 0);
      temperature_data      : in std_logic_vector(12 downto 0);
      iddt_control          : out std_logic_vector(2 downto 0);
      iddt_data             : in std_logic_vector(12 downto 0);
      slack_control         : out std_logic_vector(2 downto 0);
      slack_data            : in std_logic_vector(31 downto 0);
      voltage_control       : out std_logic_vector(2 downto 0);
      voltage_data          : in std_logic_vector(31 downto 0)
    );
end component;

	  constant clk_period : time := 10 ns;
	  constant tck_period : time := 35 ns;
    constant HALF_SEPARATOR : time := 2*tck_period;
    constant FULL_SEPARATOR : time := 8*tck_period;

	  signal reset, not_reset, clk: std_logic :='0';

    signal TCK, RST, SEL, SI, SE, UE, CE, SO, toF, toC : std_logic := '0';

    -- GPIO
    signal PE_0_GPIO_out : std_logic_vector(15 downto 0);
    signal PE_0_GPIO_in : std_logic_vector(21 downto 0) := (others => '1');
    signal uart_write_0,  uart_write_1, uart_write_2, uart_write_3: std_logic;
    signal uart_read_0,   uart_read_1,  uart_read_2,  uart_read_3: std_logic;

    signal temperature_control   : std_logic_vector(2 downto 0);
    signal temperature_data      : std_logic_vector(12 downto 0);
    signal iddt_control          : std_logic_vector(2 downto 0);
    signal iddt_data             : std_logic_vector(12 downto 0);
    signal slack_control         : std_logic_vector(2 downto 0);
    signal slack_data            : std_logic_vector(31 downto 0);
    signal voltage_control       : std_logic_vector(2 downto 0);
    signal voltage_data          : std_logic_vector(31 downto 0);

  signal current_test : string(1 to 16);
  signal RAM_readout: std_logic_vector(RAMDataSize-1 downto 0);
  signal r0_sta_value : std_logic_vector (0 to 24);
  signal slack_value : std_logic_vector (0 to 31);
  signal temp_value : std_logic_vector (0 to 31);
  signal volt_value : std_logic_vector (0 to 31);
  shared variable pre_shift, post_shift: std_logic_vector(0 to 127);
  shared variable pre_shift_len, post_shift_len : natural;
begin

    -- instantiating the top module for the network
    NoC_top: network_2x2_with_PE generic map (DATA_WIDTH  => 32, DATA_WIDTH_LV => 11)
    port map (reset, clk,
                TCK, RST, SEL, SI, SE, UE, CE, SO, toF, toC,
              PE_0_GPIO_out, PE_0_GPIO_in,
              uart_write_0, uart_read_0,
              uart_write_1, uart_read_1,
              uart_write_2, uart_read_2,
              uart_write_3, uart_read_3,

              temperature_control, temperature_data,
              iddt_control, iddt_data,
              slack_control, slack_data,
              voltage_control, voltage_data
             );

    -- Added for IJTAG

    not_reset <= not reset;

  clk_process :process
  begin
      clk <= '0';
      wait for clk_period/2;
      clk <= '1';
      wait for clk_period/2;
  end process;

  ijtag_shift_proc: process


  variable read_out_data: std_logic_vector(RAMDataSize-1 downto 0);

    variable I, J: integer := 0;
    variable stuck_at: std_logic_vector (1 downto 0) := (others => '0');
    variable address_fifo: std_logic_vector (5 downto 0) := (others => '0');

    variable address_arbiter_out: std_logic_vector (4 downto 0) := (others => '0');
    variable address_arbiter_in: std_logic_vector (4 downto 0) := (others => '0');
    variable address_arbiter_logic: std_logic_vector (8 downto 0) := (others => '0');
    variable address_lbdr: std_logic_vector (6 downto 0) := (others => '0');

       -- Generate a number of TCK ticks
    procedure tck_tick (number_of_tick : in positive) is
    begin
      for i in 1 to number_of_tick loop
        TCK <= '0';
        wait for TCK_period/2;
        TCK <= '1';
        wait for TCK_period/2;
      end loop;
    end procedure tck_tick;

    procedure tck_halftick_high is
    begin
      TCK <= '1';
      wait for TCK_period/2;
    end procedure tck_halftick_high;

    procedure tck_halftick_low is
    begin
      TCK <= '0';
      wait for TCK_period/2;
    end procedure tck_halftick_low;

     -- Shifts in specified data (Capture -> Shift -> Update)
    procedure shift_data (data : in std_logic_vector) is
    begin
       -- Capture phase
      CE <= '1';
      tck_tick(1);
      CE <= '0';
        -- Shift phase
      SE <= '1';

      if pre_shift_len > 0 then
        for i in 0 to pre_shift_len-1 loop
           SI <= pre_shift(i);
           tck_tick(1);
        end loop;
      end if ;

      for i in data'range loop
         SI <= data(i);
         tck_tick(1);
      end loop;

      if post_shift_len > 0 then
        for i in 0 to post_shift_len-1 loop
           SI <= post_shift(i);
           tck_tick(1);
        end loop;
      end if ;
      SE <= '0';
      -- Update phase
      tck_halftick_low;
      UE <= '1';
      tck_halftick_high;
      tck_halftick_low;
      UE <= '0';
      tck_halftick_high;
    end procedure shift_data;

     -- Shifts in specified data (Capture -> Shift -> Update)
    procedure shift_data_with_readout (data : in std_logic_vector; capture_data : out std_logic_vector) is
    begin
        --Capture phase
      CE <= '1';
      tck_tick(1);
      CE <= '0';
         --Shift phase
      SE <= '1';

      if pre_shift_len > 0 then
        for i in 0 to pre_shift_len-1 loop
           SI <= pre_shift(i);
           tck_tick(1);
        end loop;
      end if ;

      for i in data'range loop
         SI <= data(i);
         capture_data(i) := SO;
         tck_tick(1);
      end loop;

      if post_shift_len > 0 then
        for i in 0 to post_shift_len-1 loop
           SI <= post_shift(i);
           tck_tick(1);
        end loop;
      end if ;
      SE <= '0';
      -- Update phase
      --tck_tick(1);
      tck_halftick_low;
      UE <= '1';
      tck_halftick_high;
      tck_halftick_low;
      UE <= '0';
      tck_halftick_high;
    end procedure shift_data_with_readout;

          -- Returns all zeroes std_logic_vector of specified size
    function all_zeroes (number_of_zeroes : in positive) return std_logic_vector is
      variable zero_array : std_logic_vector(0 to number_of_zeroes-1);
    begin
      for i in zero_array'range loop
       zero_array(i) := '0';
      end loop;
      return zero_array;
    end function all_zeroes;

          -- Returns all ones std_logic_vector of specified size
    function all_ones (number_of_ones : in positive) return std_logic_vector is
      variable ones_array : std_logic_vector(0 to number_of_ones-1);
    begin
      for i in ones_array'range loop
       ones_array(i) := '1';
      end loop;
      return ones_array;
    end function all_ones;

    function reverse_vector (a: in std_logic_vector) return std_logic_vector is
      variable result: std_logic_vector(a'RANGE);
      alias aa: std_logic_vector(a'REVERSE_RANGE) is a;
  begin
      for i in aa'RANGE loop
        result(i) := aa(i);
      end loop;
      return result;
  end;

    procedure set_ram_address (address : in std_logic_vector(RAMAddrSize-1 downto 0); autoinc : in boolean; write_en : in boolean) is
      -- This function should be called in simulation when sib_mem is already opened, but sib_addr and sib_data are still closed
      -- After shifting in the provided bit vector, address sib is closed and data sib is opened
      constant open_mem_close_addr_sibs : std_logic_vector := "10";
      constant open_sib_data : std_logic := '1';
      variable autoincrement_bit : std_logic;
      variable writeen_bit : std_logic;
      variable bitstream_vector : std_logic_vector(0 to RAMAddrSize+4);
    begin
      if autoinc then
         autoincrement_bit := '1';
      else
         autoincrement_bit := '0';
      end if;
      if write_en then
         writeen_bit := '1';
      else
         writeen_bit := '0';
      end if;

      shift_data("11"&"0"); -- open sib_mem and sib_addr and close sib_data

      bitstream_vector(0 to 1) := open_mem_close_addr_sibs;
      bitstream_vector(2 to RAMAddrSize+1) := reverse_vector(address);
      bitstream_vector(RAMAddrSize+2) := autoincrement_bit;
      bitstream_vector(RAMAddrSize+3) := writeen_bit;
      bitstream_vector(RAMAddrSize+4) := open_sib_data;

      shift_data(bitstream_vector);
    end procedure set_ram_address;

    procedure get_set_data (write_data: in std_logic_vector (RAMDataSize-1 downto 0); read_data: out std_logic_vector (RAMDataSize-1 downto 0); leave_data_sib_open: in boolean) is
      -- This function should be called in simulation when sib_mem and sib_data is opened, but sib_addr is closed.
      constant open_mem_close_addr_sibs : std_logic_vector := "10";
      variable leavedatasibopen_bit : std_logic;
      variable read_data_vector : std_logic_vector (RAMDataSize-1 downto 0) := (others => '0');
      variable bitstream_vector : std_logic_vector (0 to RAMDataSize+2);
      variable readout_vector : std_logic_vector (0 to RAMDataSize+2);
    begin
      if leave_data_sib_open then
         leavedatasibopen_bit := '1';
      else
         leavedatasibopen_bit := '0';
      end if;

      tck_tick(3); --otherwise previous data can be captured

      bitstream_vector(0 to 1) := open_mem_close_addr_sibs;
      bitstream_vector(2) := leavedatasibopen_bit;
      bitstream_vector(3 to RAMDataSize+2) := reverse_vector(write_data);

      shift_data_with_readout(bitstream_vector, readout_vector);

      read_data := reverse_vector(readout_vector(3 to RAMDataSize+2));

    end procedure get_set_data;



    procedure test_ram_access is
    begin
      -- Now SIB_MEM open, SIB_ADDR closed, SIB_DATA closed
      current_test <= "ram0_addr_003   ";
      set_ram_address(X"003", true, true); -- Set WORD address to 0x003, autoincrement on, RAM write on
      -- Now SIB_MEM open, SIB_ADDR closed, SIB_DATA open
      current_test <= "ram0_write_to_3 ";
      get_set_data(X"0AA0F0F0", read_out_data, true); -- Shift in some data to write to address 0x003, increment address and leave SIB_DATA open
      -- Now SIB_MEM open, SIB_ADDR closed, SIB_DATA open
      current_test <= "ram0_write_to_4 ";
      get_set_data(X"0BB0FF00", read_out_data, true); -- Shift in some data to write to address 0x004, increment address and leave SIB_DATA open
      -- Now SIB_MEM open, SIB_ADDR closed, SIB_DATA open
      current_test <= "ram0_write_to_5C";
      get_set_data(X"0CC0F00F", read_out_data, false); -- Shift in some data to write to address 0x005, increment address and close SIB_DATA
      -- Now SIB_MEM open, SIB_ADDR closed, SIB_DATA closed

      current_test <= "ram0_addr_033   ";
      set_ram_address(X"033", true, true); -- Set WORD address to 0x033, autoincrement on, RAM write on
      -- Now SIB_MEM open, SIB_ADDR closed, SIB_DATA open
      current_test <= "ram0_write_to_33";
      get_set_data(X"0000F0F0", read_out_data, true); -- Shift in some data to write to address 0x033, increment address and leave SIB_DATA open
      -- Now SIB_MEM open, SIB_ADDR closed, SIB_DATA open
      current_test <= "ram0_write_to34C";
      get_set_data(X"0000FF00", read_out_data, false); -- Shift in some data to write to address 0x034, increment address and close SIB_DATA
      -- Now SIB_MEM open, SIB_ADDR closed, SIB_DATA closed

      RAM_readout <= (others => '0');
      current_test <= "ram0_addr_003   ";
      set_ram_address(X"003", true, false); -- Set WORD address to 0x003, autoincrement off, RAM write off
      -- Now SIB_MEM open, SIB_ADDR closed, SIB_DATA open
      current_test <= "ram0_read_003   ";
      get_set_data(X"00000000", read_out_data, true); -- Shift in some data (no write) and leave SIB_DATA open, possible to read out data from address 0x003
      -- Now SIB_MEM open, SIB_ADDR closed, SIB_DATA open
      current_test <= "ram0_read_004   ";
      get_set_data(X"00000000", read_out_data, false); -- Shift in some data (no write) and close SIB_DATA, possible to read out data from address 0x004
      -- Now SIB_MEM open, SIB_ADDR closed, SIB_DATA closed

      RAM_readout <= read_out_data; -- put data from word address 0x004

      current_test <= "close_sib_mem   ";
      shift_data("000"); -- close all but sib_ram: sib_noc & sib_sens & 3xsib_mem + opened sib_mem
      tck_tick(4);
    end procedure test_ram_access;

    variable r0_sta_value_var : std_logic_vector (0 to 24);
    variable slack_value_var : std_logic_vector (0 to 31);
    variable temp_value_var : std_logic_vector (0 to 31);
    variable volt_value_var : std_logic_vector (0 to 31);
  begin

--    the order of bits in each sib is: SXCF where S is opening bit!
--    to open sib 3 we need to shift the following: "0001"&"0000"&"0000"&"0000"&"0000"
--      * note that the shifting order is oposite!

--   Organization of IJTAG network (top level):
--            .----------.   .-----------.   .----------.
--     SI ----| sib_ram  |---| sib_sens  |---| sib_noc  |-- SO
--            '----------'   '-----------'   '----------'
--              |       |_________________________________________________.
--              |                                                         |
--              | .-----------. .-----------. .-----------. .-----------. |
--              '-| sib_ram_0 |-| sib_ram_1 |-| sib_ram_2 |-| sib_ram_3 |-'
--                '-----------' '-----------' '-----------' '-----------'
--          .-------.
--  SI -----|sib_mem|-- SO
--          '-------'
--            |    |_________________________________________________.
--            |                                                      |
--            |  .----------.                      .------------.    |
--            '--| sib_data |--------------------->| sib_addr   |----'
--               '----------'                      '------------'
--                |      |_____________               |      |______________
--                |     _____________  |              |   ______   _______  |
--                '--->|   data      |-'              '->|we,inc|-|address|-'
--                     '-------------'                   '------' '-------'
-- Auto increment bit is MSb in Address shift register
--            .-----------.
--     SI ----| sib_sens  |---------------------------------------------- SO
--            '-----------'
--              |       |_____________________________________________.
--              |                                                     |
--              | .----------. .----------. .----------. .----------. |
--              '-| sib_temp |-| sib_iddt |-| sib_slck |-| sib_volt |-'
--                '----------' '----------' '----------' '----------'
--            .-----------.
--     SI ----| sib_noc   |---------------------------------------------- SO
--            '-----------'
--              |       |_________________________________.
--              |                                         |
--              | .-------. .-------. .-------. .-------. |
--              '-| sib_0 |-| sib_1 |-| sib_2 |-| sib_3 |-'
--                '-------' '-------' '-------' '-------'
--                                               |    |_________________________________________.
--                                               |                                              |
--                                               |  .----------.              .------------.    |
--                                               '--| sib3 inj |------------->|sib3 status |----'
--                                                  '----------'              '------------'
--                                                   |      |_____________       |      |_____________
--                                                   |     _____________  |      |     _____________  |
--                                                   '--->|injection reg|-'      '--->|async adapter|-'
--                                                        '-------------'             '-------------'


    -- Reset iJTAG chain and Instruments
    RST <= '1';
    wait for tck_period;
    RST <= '0';
    SEL <= '1';
    tck_tick(4);
    reset <= '1';

-- RAM access instrument test

   reset <= '0';

   current_test <= "open_sib_ram    ";
   shift_data(fcXN&fcXN&fcXS); -- open sib_ram

   -- Test mem0
   current_test <= "open_sib_ram0   ";
   pre_shift(0 to 14) := fcXN&fcXN&fcXS&"0"&"0"&"0";
   pre_shift_len := 15;
   post_shift_len := 0;

   shift_data("1"); -- open sib_ram and sib_ram0: sib_noc & sib_sens & sib_ram & 3xsib_mem
   tck_tick(4);
   test_ram_access;

   -- Test mem1
   current_test <= "open_sib_ram1   ";
   pre_shift(0 to 13) := fcXN&fcXN&fcXS&"0"&"0";
   pre_shift_len := 14;
   post_shift(0 to 0) := "0";
   post_shift_len := 1;

   shift_data("1"); -- open sib_ram and sib_ram_1: sib_noc & sib_sens & sib_ram & 4xsib_mem
   tck_tick(4);
   test_ram_access;

   -- Test mem2
   current_test <= "open_sib_ram2   ";
   pre_shift(0 to 12) := fcXN&fcXN&fcXS&"0";
   pre_shift_len := 13;
   post_shift(0 to 1) := "00";
   post_shift_len := 2;

   shift_data("1"); -- open sib_ram and sib_ram_2: sib_noc & sib_sens & sib_ram & 4xsib_mem
   tck_tick(4);
   test_ram_access;

   -- Test mem2
   current_test <= "open_sib_ram3   ";
   pre_shift(0 to 11) := fcXN&fcXN&fcXS;
   pre_shift_len := 12;
   post_shift(0 to 2) := "000";
   post_shift_len := 3;

   shift_data("1"); -- open sib_ram and sib_ram_3: sib_noc & sib_sens & sib_ram & 4xsib_mem
   tck_tick(4);
   test_ram_access;

   current_test <= "close_sib_ram   ";
   pre_shift_len := 0;
   post_shift_len := 0;
   shift_data(fcXN&fcXN&fcXN&"0"&"0"&"0"&"0"); -- close all sibs

   -- Release chip reset
   reset <= '1';

   wait for 10us;

-- Sensors

    --temperature_data(12 downto 1) <= "000000000000";
    --temperature_data(0) <= '0';

    --current_test <= "open_sib_sens   ";
    --pre_shift_len := 0;
    --post_shift_len := 0;
    --shift_data(fcXN&fcXS&fcXN); -- open sib_sens

-- Temperature monitor test

    --current_test <= "open_sib_temp   ";
    --pre_shift(0 to 23) := fcXN&fcXS&fcXN&fcXN&fcXN&fcXS; -- (top)noc, (top)sens, volt, slack, iddt, sib_temp
    --pre_shift_len := 24;
    --post_shift(0 to 3) := fcXN; --(top)mem
    --post_shift_len := 4;

    --shift_data(""); --open sib_temp

    --current_test <= "shift_temp_setup";
    --shift_data("001000000000"&"010000000000"&"0"&"1"&"1"&"01111"); -- shift in threshold H without update

    --tck_tick(4);

    --current_test <= "temp 1          ";
    --temperature_data(12 downto 1) <= "000000000011";
    --tck_tick(1);
    --temperature_data(0) <= '1';
    --tck_tick(1);
    --temperature_data(0) <= '0';

    --tck_tick(4);

    --current_test <= "temp 2          ";
    --temperature_data(12 downto 1) <= "000000000100";
    --tck_tick(1);
    --temperature_data(0) <= '1';
    --tck_tick(1);
    --temperature_data(0) <= '0';

    --tck_tick(4);

    --current_test <= "temp 3          ";
    --temperature_data(12 downto 1) <= "000000001100";
    --tck_tick(1);
    --temperature_data(0) <= '1';
    --tck_tick(1);
    --temperature_data(0) <= '0';

    --tck_tick(4);

    --current_test <= "shift_temp_setup";
    --shift_data("001000000000"&"010000000000"&"0"&"0"&"1"&"01011"); -- shift in threshold H without update

    --tck_tick(10);

    --current_test <= "close_sib_temp  ";
    --pre_shift(0 to 23) := fcXN&fcXS&fcXN&fcXN&fcXN&fcXN; -- (top)noc, (top)sens, volt, slack, iddt, temp
    --pre_shift_len := 24;
    --post_shift(0 to 3) := fcXN; --(top)mem
    --post_shift_len := 4;

    ----shift_data(all_zeroes(32));
    --shift_data_with_readout(all_zeroes(32), temp_value_var);
    --temp_value <= reverse_vector(temp_value_var);

---- IDDt monitor test

--    current_test <= "open_sib_iddt   ";
--    pre_shift(0 to 19) := fcXN&fcXS&fcXN&fcXN&fcXS; -- (top)noc, (top)sens, volt, slack, iddt
--    pre_shift_len := 20;
--    post_shift(0 to 7) := fcXN&fcXN; -- temp, (top)mem
--    post_shift_len := 8;

--    shift_data(""); --open sib_temp


--    current_test <= "close_sib_iddt  ";
--    pre_shift(0 to 19) := fcXN&fcXS&fcXN&fcXN&fcXN; -- (top)noc, (top)sens, volt, slack, iddt
--    pre_shift_len := 20;
--    post_shift(0 to 7) := fcXN&fcXN; -- temp, (top)mem
--    post_shift_len := 8;

--    shift_data(all_zeroes(32));

-- Slack monitor test

    --current_test <= "open_sib_slack  ";
    --pre_shift(0 to 15) := fcXN&fcXS&fcXN&fcXS; -- (top)noc, (top)sens, volt, slack
    --pre_shift_len := 16;
    --post_shift(0 to 11) := fcXN&fcXN&fcXN; -- iddt, temp, (top)mem
    --post_shift_len := 12;

    --shift_data(""); --open sib_temp

    --current_test <= "Slack           ";
    --shift_data("11100"&"00000"&"0"&"1"&"1"&"0000000000000001111"); -- shift in threshold H without update
    --tck_tick(4);

    --slack_data <= "00101010101010101010101010101010";
    --tck_tick(10);
    --slack_data <= "10101010101010101010101010100101";
    --tck_tick(4);

    --current_test <= "close_sib_slack ";
    --pre_shift(0 to 15) := fcXN&fcXS&fcXN&fcXN; -- (top)noc, (top)sens, volt, slack
    --pre_shift_len := 16;
    --post_shift(0 to 11) := fcXN&fcXN&fcXN; -- iddt, temp, (top)mem
    --post_shift_len := 12;

    --shift_data_with_readout(all_zeroes(32), slack_value_var);
    --slack_value <= reverse_vector(slack_value_var);
    --shift_data(all_zeroes(32));

-- Voltage monitor test

    --voltage_data <= "00000000000000000000000000000000";

    --current_test <= "open_sib_volt   ";
    --pre_shift(0 to 11) := fcXN&fcXS&fcXS; -- (top)noc, (top)sens, volt
    --pre_shift_len := 12;
    --post_shift(0 to 15) := fcXN&fcXN&fcXN&fcXN; -- slack, iddt, temp, (top)mem
    --post_shift_len := 16;

    --shift_data(""); --open sib_temp

    --current_test <= "Voltage         ";
    --shift_data("00001"&"11100"&"1"&"1"&"1"&"0000000000000001111"); -- shift in threshold H without update

    --voltage_data <= "00000000000000000000000000000000";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000000000000001";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000000000000011";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000000000000111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000000000001111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000000000011111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000000000111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000000001111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000000011111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000000111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000001111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000011111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000000111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000001111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000011111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000000111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000001111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000011111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000000111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000001111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000011111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000000111111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000001111111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000011111111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000000111111111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000001111111111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000011111111111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00000111111111111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00001111111111111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00011111111111111111111111111111";
    --tck_tick(1);
    --voltage_data <= "00111111111111111111111111111111";
    --tck_tick(1);
    --voltage_data <= "01111111111111111111111111111111";
    --tck_tick(1);
    --voltage_data <= "11111111111111111111111111111111";
    --tck_tick(10);

    --shift_data("11100"&"00001"&"0"&"1"&"1"&"0000000000000001111"); -- shift in threshold H without update
    --tck_tick(10);

    --voltage_data <= "00000000000000000000000011111111";
    --tck_tick(10);

    --current_test <= "close_sib_volt  ";
    --pre_shift(0 to 11) := fcXN&fcXS&fcXN; -- (top)noc, (top)sens, volt
    --pre_shift_len := 12;
    --post_shift(0 to 15) := fcXN&fcXN&fcXN&fcXN; -- slack, iddt, temp, (top)mem
    --post_shift_len := 16;

    ----shift_data(all_zeroes(32));
    --shift_data_with_readout(all_zeroes(32), volt_value_var);
    --volt_value <= reverse_vector(volt_value_var);

    --current_test <= "close_sib_sens  ";
    --pre_shift_len := 0;
    --post_shift_len := 0;
    --shift_data(fcXN&fcXN&fcXN&fcXN&fcXN&fcXN&fcXN); -- close all sibs

-- Router SIBs

    current_test <= "open_sib_noc    ";
    pre_shift_len := 0;
    post_shift_len := 0;
    shift_data(fcXS&fcXN&fcXN); -- open sib_noc

    --Router 0
    current_test <= "open_sib_r0     ";
    pre_shift(0 to 19) := fcXS&fcXN&fcXN&fcXN&fcXS; -- (top)noc, r3, r2, r1, r0
    pre_shift_len := 20;
    post_shift(0 to 7) := fcXN&fcXN; -- (top)sens, (top)mem
    post_shift_len := 8;

    shift_data(""); --open sib_r0

    --Router 0 injection
    current_test <= "open_sib_r0_inj ";
    pre_shift(0 to 27) := fcXS&fcXN&fcXN&fcXN&fcXS&fcXN&fcXS; -- (top)noc, r3, r2, r1, r0, r0_sta, r0_inj
    pre_shift_len := 28;
    post_shift(0 to 7) := fcXN&fcXN; -- (top)sens, (top)mem
    post_shift_len := 8;

    shift_data(""); --open sib_r0_inj

    current_test <= "r0_inj_arb_out  ";
    --shift_data(all_zeroes(130));
    shift_data("000000000"&   "0000001"&"0000001"&"0000001"&"0000001"&"0000001"&   "0000000"&"0000000"&"0000000"&"0000000"&"0000000"&   "000000000"&"000000000"&"000000000"&   "00000000"&"00000000"&"00000000");


    current_test <= "close_sib_r0_inj";
    pre_shift(0 to 27) := fcXS&fcXN&fcXN&fcXN&fcXS&fcXN&fcXN; -- (top)noc, r3, r2, r1, r0, r0_sta, r0_inj
    pre_shift_len := 28;
    post_shift(0 to 7) := fcXN&fcXN; -- (top)sens, (top)mem
    post_shift_len := 8;

    shift_data(all_zeroes(130));

    --Router 0 status
    current_test <= "open_sib_r0_sta ";
    pre_shift(0 to 23) := fcXS&fcXN&fcXN&fcXN&fcXS&fcXS; -- (top)noc, r3, r2, r1, r0, r0_sta
    pre_shift_len := 24;
    post_shift(0 to 11) := fcXN&fcXN&fcXN; -- r0_inj, (top)sens, (top)mem
    post_shift_len := 12;

    shift_data(""); --open sib_r0_sta

    current_test <= "r0_sta_readout  ";
    shift_data_with_readout(all_zeroes(25), r0_sta_value_var);
    r0_sta_value <= reverse_vector(r0_sta_value_var);
    --shift_data(all_zeroes(25));


    current_test <= "close_sib_r0_sta";
    pre_shift(0 to 23) := fcXS&fcXN&fcXN&fcXN&fcXS&fcXN; -- (top)noc, r3, r2, r1, r0, r0_sta
    pre_shift_len := 24;
    post_shift(0 to 11) := fcXN&fcXN&fcXN; -- r0_inj, (top)sens, (top)mem
    post_shift_len := 12;

    shift_data("11111"&all_zeroes(20));

    current_test <= "close_sib_r0    ";
    pre_shift(0 to 19) := fcXS&fcXN&fcXN&fcXN&fcXN; -- (top)noc, r3, r2, r1, r0
    pre_shift_len := 20;
    post_shift(0 to 7) := fcXN&fcXN; -- (top)sens, (top)mem
    post_shift_len := 8;

    shift_data(fcXN&fcXN); -- inj and status sibs of r0






    ----Router 1
    --current_test <= "open_sib_r1     ";
    --pre_shift(0 to 15) := fcXS&fcXN&fcXN&fcXS; -- (top)noc, r3, r2, r1
    --pre_shift_len := 16;
    --post_shift(0 to 11) := fcXN&fcXN&fcXN; -- r0, (top)sens, (top)mem
    --post_shift_len := 12;

    --shift_data(""); --open sib_r1

    ----Router 1 injection
    --current_test <= "open_sib_r1_inj ";
    --pre_shift(0 to 23) := fcXS&fcXN&fcXN&fcXS&fcXN&fcXS; -- (top)noc, r3, r2, r1, r1_sta, r1_inj
    --pre_shift_len := 24;
    --post_shift(0 to 11) := fcXN&fcXN&fcXN; -- r0, (top)sens, (top)mem
    --post_shift_len := 12;

    --shift_data(""); --open sib_r1_inj

    --current_test <= "r1_inj_arb_out  ";
    --shift_data(all_zeroes(130));
    ----shift_data("000000000"&   "0000001"&"0000001"&"0000001"&"0000001"&"0000001"&   "0000000"&"0000000"&"0000000"&"0000000"&"0000000"&   "000000000"&"000000000"&"000000000"&   "00000000"&"00000000"&"00000000");


    --current_test <= "close_sib_r1_inj";
    --pre_shift(0 to 23) := fcXS&fcXN&fcXN&fcXS&fcXN&fcXN; -- (top)noc, r3, r2, r1, r1_sta, r1_inj
    --pre_shift_len := 24;
    --post_shift(0 to 11) := fcXN&fcXN&fcXN; -- r0, (top)sens, (top)mem
    --post_shift_len := 12;

    --shift_data(all_zeroes(130));

    --current_test <= "close_sib_r1    ";
    --pre_shift(0 to 15) := fcXS&fcXN&fcXN&fcXN; -- (top)noc, r3, r2, r1
    --pre_shift_len := 16;
    --post_shift(0 to 11) := fcXN&fcXN&fcXN; -- r0, (top)sens, (top)mem
    --post_shift_len := 12;

    --shift_data(fcXN&fcXN); -- inj and status sibs of r1

    ----Router 2
    --current_test <= "open_sib_r2     ";
    --pre_shift(0 to 11) := fcXS&fcXN&fcXS; -- (top)noc, r3, r2
    --pre_shift_len := 12;
    --post_shift(0 to 15) := fcXN&fcXN&fcXN&fcXN; -- r1, r0, (top)sens, (top)mem
    --post_shift_len := 16;

    --shift_data(""); --open sib_r2

    ----Router 2 injection
    --current_test <= "open_sib_r2_inj ";
    --pre_shift(0 to 19) := fcXS&fcXN&fcXS&fcXN&fcXS; -- (top)noc, r3, r2, r2_sta, r2_inj
    --pre_shift_len := 20;
    --post_shift(0 to 15) := fcXN&fcXN&fcXN&fcXN; -- r1, r0, (top)sens, (top)mem
    --post_shift_len := 16;

    --shift_data(""); --open sib_r2_inj

    --current_test <= "r2_inj_arb_out  ";
    --shift_data(all_zeroes(130));
    ----shift_data("000000000"&   "0000001"&"0000001"&"0000001"&"0000001"&"0000001"&   "0000000"&"0000000"&"0000000"&"0000000"&"0000000"&   "000000000"&"000000000"&"000000000"&   "00000000"&"00000000"&"00000000");


    --current_test <= "close_sib_r2_inj";
    --pre_shift(0 to 19) := fcXS&fcXN&fcXS&fcXN&fcXN; -- (top)noc, r3, r2, r2_sta, r2_inj
    --pre_shift_len := 20;
    --post_shift(0 to 15) := fcXN&fcXN&fcXN&fcXN; -- r1, r0, (top)sens, (top)mem
    --post_shift_len := 16;

    --shift_data(all_zeroes(130));


    --current_test <= "close_sib_r2    ";
    --pre_shift(0 to 11) := fcXS&fcXN&fcXN; -- (top)noc, r3, r2
    --pre_shift_len := 12;
    --post_shift(0 to 15) := fcXN&fcXN&fcXN&fcXN; -- r1, r0, (top)sens, (top)mem
    --post_shift_len := 16;

    --shift_data(fcXN&fcXN); -- inj and status sibs of r2

    ----Router 3
    --current_test <= "open_sib_r3     ";
    --pre_shift(0 to 7) := fcXS&fcXS; -- (top)noc, r3
    --pre_shift_len := 8;
    --post_shift(0 to 19) := fcXN&fcXN&fcXN&fcXN&fcXN; -- r2, r1, r0, (top)sens, (top)mem
    --post_shift_len := 20;

    --shift_data(""); --open sib_r3

    ----Router 2 injection
    --current_test <= "open_sib_r3_inj ";
    --pre_shift(0 to 15) := fcXS&fcXS&fcXN&fcXS; -- (top)noc, r3, r3_sta, r3_inj
    --pre_shift_len := 16;
    --post_shift(0 to 19) := fcXN&fcXN&fcXN&fcXN&fcXN; -- r2, r1, r0, (top)sens, (top)mem
    --post_shift_len := 20;

    --shift_data(""); --open sib_r3_inj

    --current_test <= "r3_inj_arb_out  ";
    --shift_data(all_zeroes(130));
    ----shift_data("000000000"&   "0000001"&"0000001"&"0000001"&"0000001"&"0000001"&   "0000000"&"0000000"&"0000000"&"0000000"&"0000000"&   "000000000"&"000000000"&"000000000"&   "00000000"&"00000000"&"00000000");


    --current_test <= "close_sib_r3_inj";
    --pre_shift(0 to 15) := fcXS&fcXS&fcXN&fcXN; -- (top)noc, r3, r3_sta, r3_inj
    --pre_shift_len := 16;
    --post_shift(0 to 19) := fcXN&fcXN&fcXN&fcXN&fcXN; -- r2, r1, r0, (top)sens, (top)mem
    --post_shift_len := 20;

    --shift_data(all_zeroes(130));

    --current_test <= "close_sib_r3    ";
    --pre_shift(0 to 7) := fcXS&fcXN; -- (top)noc, r3
    --pre_shift_len := 8;
    --post_shift(0 to 19) := fcXN&fcXN&fcXN&fcXN&fcXN; -- r2, r1, r0, (top)sens, (top)mem
    --post_shift_len := 20;

    --shift_data(fcXN&fcXN); -- inj and status sibs of r3




    current_test <= "close_sib_noc   ";
    pre_shift_len := 0;
    post_shift_len := 0;
    shift_data(fcXN&fcXN&fcXN&fcXN&fcXN&fcXN&fcXN); -- close all sibs

    wait;

end process;

end behavior;
