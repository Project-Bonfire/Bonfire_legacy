--Copyright (C) 2016 Siavoosh Payandeh Azad
------------------------------------------------------------
-- This file is automatically generated!
-- Here are the parameters:
-- 	 network size x: 2
-- 	 network size y: 2
-- 	 Data width: 32
-- 	 Parity: False
------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ieee.numeric_std.ALL; 
use work.component_pack.all;
use ieee.std_logic_misc.all;

entity network_2x2 is
 generic (DATA_WIDTH: integer := 32; DATA_WIDTH_LV: integer := 11);
port (reset: in  std_logic; 
	clk: in  std_logic; 
	--------------
	--------------
	RX_L_0: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_0, valid_out_L_0: out std_logic;
	credit_in_L_0, valid_in_L_0: in std_logic;
	TX_L_0: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_1: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_1, valid_out_L_1: out std_logic;
	credit_in_L_1, valid_in_L_1: in std_logic;
	TX_L_1: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_2: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_2, valid_out_L_2: out std_logic;
	credit_in_L_2, valid_in_L_2: in std_logic;
	TX_L_2: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
	RX_L_3: in std_logic_vector (DATA_WIDTH-1 downto 0);
	credit_out_L_3, valid_out_L_3: out std_logic;
	credit_in_L_3, valid_in_L_3: in std_logic;
	TX_L_3: out std_logic_vector (DATA_WIDTH-1 downto 0);
	--------------
    link_faults_0: out std_logic_vector(4 downto 0);
    turn_faults_0: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_0: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_0: in  std_logic_vector(3 downto 0);
    Reconfig_command_0 : in std_logic;

	--------------
    link_faults_1: out std_logic_vector(4 downto 0);
    turn_faults_1: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_1: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_1: in  std_logic_vector(3 downto 0);
    Reconfig_command_1 : in std_logic;

	--------------
    link_faults_2: out std_logic_vector(4 downto 0);
    turn_faults_2: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_2: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_2: in  std_logic_vector(3 downto 0);
    Reconfig_command_2 : in std_logic;

	--------------
    link_faults_3: out std_logic_vector(4 downto 0);
    turn_faults_3: out std_logic_vector(19 downto 0);
    Rxy_reconf_PE_3: in  std_logic_vector(7 downto 0);
    Cx_reconf_PE_3: in  std_logic_vector(3 downto 0);
    Reconfig_command_3 : in std_logic;

    --------------
    -- IJTAG network for fault injection and checker status monitoring
    TCK         : in std_logic;
    RST         : in std_logic;
    SEL         : in std_logic;
    SI          : in std_logic;
    SE          : in std_logic;
    UE          : in std_logic;
    CE          : in std_logic;
    SO          : out std_logic;
    toF         : out std_logic;
    toC         : out std_logic
    ); 
end network_2x2; 


architecture behavior of network_2x2 is


-- For IJAG

component SIB_mux_pre_FCX_SELgate is
    Port ( -- Scan Interface  client --------------
           SI : in STD_LOGIC; -- ScanInPort 
           CE : in STD_LOGIC; -- CaptureEnPort
           SE : in STD_LOGIC; -- ShiftEnPort
           UE : in STD_LOGIC; -- UpdateEnPort
           SEL : in STD_LOGIC; -- SelectPort
           RST : in STD_LOGIC; -- ResetPort
           TCK : in STD_LOGIC; -- TCKPort
           SO : out STD_LOGIC; -- ScanOutPort
           toF : out STD_LOGIC; -- To F flag of the upper hierarchical level
           toC : out STD_LOGIC; -- To C flag of the upper hierarchical level
       -- Scan Interface  host ----------------
           fromSO : in  STD_LOGIC; -- ScanInPort
           toCE : out  STD_LOGIC; -- ToCaptureEnPort
           toSE : out  STD_LOGIC; -- ToShiftEnPort
           toUE : out  STD_LOGIC; -- ToUpdateEnPort
           toSEL : out  STD_LOGIC; -- ToSelectPort
           toRST : out  STD_LOGIC; -- ToResetPort
           toTCK : out  STD_LOGIC; -- ToTCKPort
           toSI : out  STD_LOGIC; -- ScanOutPort
           fromF : in STD_LOGIC; -- From an OR of all F flags in the underlying network segment
           fromC : in STD_LOGIC);  -- From an AND of all C flags in the underlying network segment
end component;

component AsyncDataRegisterAdapter is
 Generic ( Size : positive);
    Port ( -- Scan Interface scan_client ----------
           SI : in STD_LOGIC; -- ScanInPort 
           SO : out STD_LOGIC; -- ScanOutPort
           SEL : in STD_LOGIC; -- SelectPort
           ----------------------------------------     
           SE : in STD_LOGIC; -- ShiftEnPort
           CE : in STD_LOGIC; -- CaptureEnPort
           UE : in STD_LOGIC; -- UpdateEnPort
           RST : in STD_LOGIC; -- ResetPort
           TCK : in STD_LOGIC; -- TCKPort
              -- Data interface
           DI : in STD_LOGIC_VECTOR (Size-1 downto 0);
           DO : out STD_LOGIC_VECTOR (Size-1 downto 0));
end component;


-- generating bulk signals. not all of them are used in the design...
	signal credit_out_N_0, credit_out_E_0, credit_out_W_0, credit_out_S_0: std_logic;
	signal credit_out_N_1, credit_out_E_1, credit_out_W_1, credit_out_S_1: std_logic;
	signal credit_out_N_2, credit_out_E_2, credit_out_W_2, credit_out_S_2: std_logic;
	signal credit_out_N_3, credit_out_E_3, credit_out_W_3, credit_out_S_3: std_logic;

	signal credit_in_N_0, credit_in_E_0, credit_in_W_0, credit_in_S_0: std_logic;
	signal credit_in_N_1, credit_in_E_1, credit_in_W_1, credit_in_S_1: std_logic;
	signal credit_in_N_2, credit_in_E_2, credit_in_W_2, credit_in_S_2: std_logic;
	signal credit_in_N_3, credit_in_E_3, credit_in_W_3, credit_in_S_3: std_logic;

	signal RX_N_0, RX_E_0, RX_W_0, RX_S_0 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_1, RX_E_1, RX_W_1, RX_S_1 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_2, RX_E_2, RX_W_2, RX_S_2 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal RX_N_3, RX_E_3, RX_W_3, RX_S_3 : std_logic_vector (DATA_WIDTH-1 downto 0);

	signal valid_out_N_0, valid_out_E_0, valid_out_W_0, valid_out_S_0: std_logic;
	signal valid_out_N_1, valid_out_E_1, valid_out_W_1, valid_out_S_1: std_logic;
	signal valid_out_N_2, valid_out_E_2, valid_out_W_2, valid_out_S_2: std_logic;
	signal valid_out_N_3, valid_out_E_3, valid_out_W_3, valid_out_S_3: std_logic;

	signal valid_in_N_0, valid_in_E_0, valid_in_W_0, valid_in_S_0: std_logic;
	signal valid_in_N_1, valid_in_E_1, valid_in_W_1, valid_in_S_1: std_logic;
	signal valid_in_N_2, valid_in_E_2, valid_in_W_2, valid_in_S_2: std_logic;
	signal valid_in_N_3, valid_in_E_3, valid_in_W_3, valid_in_S_3: std_logic;

	signal TX_N_0, TX_E_0, TX_W_0, TX_S_0 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_1, TX_E_1, TX_W_1, TX_S_1 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_2, TX_E_2, TX_W_2, TX_S_2 : std_logic_vector (DATA_WIDTH-1 downto 0);
	signal TX_N_3, TX_E_3, TX_W_3, TX_S_3 : std_logic_vector (DATA_WIDTH-1 downto 0);

	signal Faulty_N_out0,Faulty_E_out0,Faulty_W_out0,Faulty_S_out0: std_logic;
	signal Faulty_N_in0,Faulty_E_in0,Faulty_W_in0,Faulty_S_in0: std_logic;
	signal Faulty_N_out1,Faulty_E_out1,Faulty_W_out1,Faulty_S_out1: std_logic;
	signal Faulty_N_in1,Faulty_E_in1,Faulty_W_in1,Faulty_S_in1: std_logic;
	signal Faulty_N_out2,Faulty_E_out2,Faulty_W_out2,Faulty_S_out2: std_logic;
	signal Faulty_N_in2,Faulty_E_in2,Faulty_W_in2,Faulty_S_in2: std_logic;
	signal Faulty_N_out3,Faulty_E_out3,Faulty_W_out3,Faulty_S_out3: std_logic;
	signal Faulty_N_in3,Faulty_E_in3,Faulty_W_in3,Faulty_S_in3: std_logic;

    -- fault injector signals
    signal TCK_0, TCK_1, TCK_2, TCK_3: std_logic;
    signal SE_0,  SE_1,  SE_2,  SE_3:  std_logic;
    signal UE_0,  UE_1,  UE_2,  UE_3:  std_logic;
    signal SI_0,  SI_1,  SI_2,  SI_3:  std_logic;
    signal SO_0,  SO_1,  SO_2,  SO_3:  std_logic;

    --------------
    -- IJTAG network signals
    signal SIB_0_toSEL,  SIB_1_toSEL,  SIB_2_toSEL,  SIB_3_toSEL  : std_logic;
    signal SIB_0_toCE,   SIB_1_toCE,   SIB_2_toCE,   SIB_3_toCE   : std_logic;
    signal SIB_0_toSE,   SIB_1_toSE,   SIB_2_toSE,   SIB_3_toSE   : std_logic;
    signal SIB_0_toUE,   SIB_1_toUE,   SIB_2_toUE,   SIB_3_toUE   : std_logic;
    signal SIB_0_toSI,   SIB_1_toSI,   SIB_2_toSI,   SIB_3_toSI   : std_logic;
    signal SIB_0_toRST,  SIB_1_toRST,  SIB_2_toRST,  SIB_3_toRST  : std_logic;
    signal SIB_0_toTCK,  SIB_1_toTCK,  SIB_2_toTCK,  SIB_3_toTCK  : std_logic;
    signal SIB_0_so,     SIB_1_so,     SIB_2_so,     SIB_3_so     : std_logic;
        
    signal SIB_0_inj_toSI,  SIB_1_inj_toSI,  SIB_2_inj_toSI,  SIB_3_inj_toSI  : std_logic;    
    signal SIB_0_inj_toTCK, SIB_1_inj_toTCK, SIB_2_inj_toTCK, SIB_3_inj_toTCK : std_logic;    
    signal SIB_0_inj_toRST, SIB_1_inj_toRST, SIB_2_inj_toRST, SIB_3_inj_toRST : std_logic;    
    signal SIB_0_inj_toSEL, SIB_1_inj_toSEL, SIB_2_inj_toSEL, SIB_3_inj_toSEL : std_logic;    
    signal SIB_0_inj_toUE,  SIB_1_inj_toUE,  SIB_2_inj_toUE,  SIB_3_inj_toUE  : std_logic;    
    signal SIB_0_inj_toSE,  SIB_1_inj_toSE,  SIB_2_inj_toSE,  SIB_3_inj_toSE  : std_logic;
    signal SIB_0_inj_toCE,  SIB_1_inj_toCE,  SIB_2_inj_toCE,  SIB_3_inj_toCE  : std_logic;
    signal SIB_0_inj_so,    SIB_1_inj_so,    SIB_2_inj_so,    SIB_3_inj_so    : std_logic;
    
    signal SIB_0_sta_toSI,  SIB_1_sta_toSI,  SIB_2_sta_toSI,  SIB_3_sta_toSI  : std_logic;    
    signal SIB_0_sta_toTCK, SIB_1_sta_toTCK, SIB_2_sta_toTCK, SIB_3_sta_toTCK : std_logic;    
    signal SIB_0_sta_toRST, SIB_1_sta_toRST, SIB_2_sta_toRST, SIB_3_sta_toRST : std_logic;    
    signal SIB_0_sta_toSEL, SIB_1_sta_toSEL, SIB_2_sta_toSEL, SIB_3_sta_toSEL : std_logic;    
    signal SIB_0_sta_toUE,  SIB_1_sta_toUE,  SIB_2_sta_toUE,  SIB_3_sta_toUE  : std_logic;    
    signal SIB_0_sta_toSE,  SIB_1_sta_toSE,  SIB_2_sta_toSE,  SIB_3_sta_toSE  : std_logic;
    signal SIB_0_sta_toCE,  SIB_1_sta_toCE,  SIB_2_sta_toCE,  SIB_3_sta_toCE  : std_logic;
    signal SIB_0_sta_so,    SIB_1_sta_so,    SIB_2_sta_so,    SIB_3_sta_so    : std_logic;

    signal SIB_main_toCE, SIB_main_toSE, SIB_main_toUE, SIB_main_toSEL, SIB_main_toRST, SIB_main_toTCK, SIB_main_toSI, toF_SIB_main, toC_SIB_main : std_logic;

    -- flags from checkers
    signal F_R0, F_R1, F_R2, F_R3 : std_logic;
    signal C_R0, C_R1, C_R2, C_R3 : std_logic;
    -- flags top level
    signal F_segtop_fromSIB_0, C_segtop_fromSIB_0 : std_logic;
    signal F_segtop_fromSIB_1, C_segtop_fromSIB_1 : std_logic;
    signal F_segtop_fromSIB_2, C_segtop_fromSIB_2 : std_logic;
    signal F_segtop_fromSIB_3, C_segtop_fromSIB_3 : std_logic;
    -- flags second level
    signal toF_SIB_0,          toF_SIB_1,          toF_SIB_2,          toF_SIB_3          : std_logic;
    signal toC_SIB_0,          toC_SIB_1,          toC_SIB_2,          toC_SIB_3          : std_logic;
    signal F_fromSIB_0_inj,    F_fromSIB_1_inj,    F_fromSIB_2_inj,    F_fromSIB_3_inj    : std_logic;
    signal C_fromSIB_0_inj,    C_fromSIB_1_inj,    C_fromSIB_2_inj,    C_fromSIB_3_inj    : std_logic;
    signal F_fromSIB_0_status, F_fromSIB_1_status, F_fromSIB_2_status, F_fromSIB_3_status : std_logic;
    signal C_fromSIB_0_status, C_fromSIB_1_status, C_fromSIB_2_status, C_fromSIB_3_status : std_logic;

    signal R0_inj_so,         R1_inj_so,         R2_inj_so,         R3_inj_so         : std_logic;
    signal R0_sta_adapter_so, R1_sta_adapter_so, R2_sta_adapter_so, R3_sta_adapter_so : std_logic;
    signal R0_sta_adapter_do, R1_sta_adapter_do, R2_sta_adapter_do, R3_sta_adapter_do : std_logic_vector(24 downto 0);
    
    signal R0_aggregated_fault_status, R1_aggregated_fault_status, R2_aggregated_fault_status, R3_aggregated_fault_status : std_logic_vector(24 downto 0);

    --------------
    -- the checker output related ports (for unclassified fault information)
    signal link_faults_async_0 : std_logic_vector(4 downto 0);
    signal turn_faults_async_0: std_logic_vector(19 downto 0);
    --------------
    signal link_faults_async_1 : std_logic_vector(4 downto 0);
    signal turn_faults_async_1: std_logic_vector(19 downto 0);
    --------------
    signal link_faults_async_2 : std_logic_vector(4 downto 0);
    signal turn_faults_async_2: std_logic_vector(19 downto 0);
    --------------
    signal link_faults_async_3 : std_logic_vector(4 downto 0);
    signal turn_faults_async_3: std_logic_vector(19 downto 0);
    --------------
--        organizaiton of the network:
--     x --------------->
--  y         ----       ----
--  |        | 0  | --- | 1  |
--  |         ----       ----
--  |          |          |
--  |         ----       ----
--  |        | 2  | --- | 3  |
--  v         ----       ----
--

--   Organization of IJTAG network (NoC part):
--            .-----------.                                    
--     SI ----| sib_main  |---------------------------------------------- SO
--            '-----------'                               
--              |       |_________________________________. 
--              |                                         | 
--              | .-------. .-------. .-------. .-------. | 
--              '-| sib_0 |-| sib_1 |-| sib_2 |-| sib_3 |-' 
--                '-------' '-------' '-------' '-------'   
--                                               |    |_________________________________________.
--                                               |                                              |
--                                               |  .----------.              .------------.    |
--                                               '--| sib3 inj |------------->|sib3 status |----'
--                                                  '----------'              '------------'
--                                                   |      |_____________       |      |_____________
--                                                   |     _____________  |      |     _____________  |
--                                                   '--->|injection reg|-'      '--->|async adapter|-'
--                                                        '-------------'             '-------------'
--
--    the order of bits in each sib is: SXCF where S is opening bit!

begin

-- IJTAG top level

SIB_main : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI  => SI,
    CE  => CE,
    SE  => SE,
    UE  => UE,
    SEL => SEL,
    RST => RST,
    TCK => TCK,
    SO  => SO,
    toF => toF,
    toC => toC,
     -- Scan Interface  host ----------------
    fromSO => SIB_3_so,
    toCE   => SIB_main_toCE,
    toSE   => SIB_main_toSE,
    toUE   => SIB_main_toUE,
    toSEL  => SIB_main_toSEL,
    toRST  => SIB_main_toRST,
    toTCK  => SIB_main_toTCK,
    toSI   => SIB_main_toSI,
    fromF  => toF_SIB_main,
    fromC  => toC_SIB_main
);

toF_SIB_main <= F_segtop_fromSIB_0 or  F_segtop_fromSIB_1 or  F_segtop_fromSIB_2 or  F_segtop_fromSIB_3;
toC_SIB_main <= C_segtop_fromSIB_0 and C_segtop_fromSIB_1 and C_segtop_fromSIB_2 and C_segtop_fromSIB_3;

-----------------------------------
------ ROUTER 0 -------------------
-----------------------------------
-- Router 0 main SIB
SIB_0 : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_main_toSI,
    CE => SIB_main_toCE,
    SE => SIB_main_toSE,
    UE => SIB_main_toUE,
    SEL => SIB_main_toSEL,
    RST => SIB_main_toRST,
    TCK => SIB_main_toTCK,
    SO => SIB_0_so,
    toF => F_segtop_fromSIB_0,
    toC => C_segtop_fromSIB_0,
     -- Scan Interface  host ----------------
    fromSO => SIB_0_sta_so,
    toCE => SIB_0_toCE,
    toSE => SIB_0_toSE,
    toUE => SIB_0_toUE,
    toSEL => SIB_0_toSEL,
    toRST => SIB_0_toRST,
    toTCK => SIB_0_toTCK,
    toSI => SIB_0_toSI,
    fromF => toF_SIB_0,
    fromC => toC_SIB_0
);

toF_SIB_0 <= F_fromSIB_0_inj or  F_fromSIB_0_status;
toC_SIB_0 <= C_fromSIB_0_inj and C_fromSIB_0_status;

-- Router 0 fault injection SIB
SIB_0_injection : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_0_toSI,
    CE => SIB_0_toCE,
    SE => SIB_0_toSE,
    UE => SIB_0_toUE,
    SEL => SIB_0_toSEL,
    RST => SIB_0_toRST,
    TCK => SIB_0_toTCK,
    SO => SIB_0_inj_so,
    toF => F_fromSIB_0_inj,
    toC => C_fromSIB_0_inj,
     -- Scan Interface  host ----------------
    fromSO => R0_inj_so,
    toCE => SIB_0_inj_toCE,
    toSE => SIB_0_inj_toSE,
    toUE => SIB_0_inj_toUE,
    toSEL => SIB_0_inj_toSEL,
    toRST => SIB_0_inj_toRST,
    toTCK => SIB_0_inj_toTCK,
    toSI => SIB_0_inj_toSI,
    fromF => '0',
    fromC => '1'
);
-- Router 0 checker status SIB
SIB_0_status : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_0_inj_so,
    CE => SIB_0_toCE,
    SE => SIB_0_toSE,
    UE => SIB_0_toUE,
    SEL => SIB_0_toSEL,
    RST => SIB_0_toRST,
    TCK => SIB_0_toTCK,
    SO => SIB_0_sta_so,
    toF => F_fromSIB_0_status,
    toC => C_fromSIB_0_status,
     -- Scan Interface  host ----------------
    fromSO => R0_sta_adapter_so,
    toCE => SIB_0_sta_toCE,
    toSE => SIB_0_sta_toSE,
    toUE => SIB_0_sta_toUE,
    toSEL => SIB_0_sta_toSEL,
    toRST => SIB_0_sta_toRST,
    toTCK => SIB_0_sta_toTCK,
    toSI => SIB_0_sta_toSI,
    fromF => F_R0,
    fromC => C_R0
);
-- Router 0 checker status IJTAG adapter
R0_status_adapter : AsyncDataRegisterAdapter
    generic map (Size => 25)
    port map (
    SI => SIB_0_sta_toSI,
    SO => R0_sta_adapter_so,
    SEL => SIB_0_sta_toSEL,
    ----------------------------------------     
    SE => SIB_0_sta_toSE,
    CE => SIB_0_sta_toCE,
    UE => SIB_0_sta_toUE,
    RST => SIB_0_sta_toRST,
    TCK => SIB_0_sta_toTCK,
      -- Data interface
    DI => R0_aggregated_fault_status,
    DO => R0_sta_adapter_do
);

R0_aggregated_fault_status <= link_faults_async_0 & turn_faults_async_0;
-----------------------------------
------ ROUTER 1 -------------------
-----------------------------------
-- Router 1 main SIB
SIB_1 : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_0_so,
    CE => SIB_main_toCE,
    SE => SIB_main_toSE,
    UE => SIB_main_toUE,
    SEL => SIB_main_toSEL,
    RST => SIB_main_toRST,
    TCK => SIB_main_toTCK,
    SO => SIB_1_so,
    toF => F_segtop_fromSIB_1,
    toC => C_segtop_fromSIB_1,
     -- Scan Interface  host ----------------
    fromSO => SIB_1_sta_so,
    toCE => SIB_1_toCE,
    toSE => SIB_1_toSE,
    toUE => SIB_1_toUE,
    toSEL => SIB_1_toSEL,
    toRST => SIB_1_toRST,
    toTCK => SIB_1_toTCK,
    toSI => SIB_1_toSI,
    fromF => toF_SIB_1,
    fromC => toC_SIB_1
);

toF_SIB_1 <= F_fromSIB_1_inj or  F_fromSIB_1_status;
toC_SIB_1 <= C_fromSIB_1_inj and C_fromSIB_1_status;

-- Router 1 fault injection SIB
SIB_1_injection : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_1_toSI,
    CE => SIB_1_toCE,
    SE => SIB_1_toSE,
    UE => SIB_1_toUE,
    SEL => SIB_1_toSEL,
    RST => SIB_1_toRST,
    TCK => SIB_1_toTCK,
    SO => SIB_1_inj_so,
    toF => F_fromSIB_1_inj,
    toC => C_fromSIB_1_inj,
     -- Scan Interface  host ----------------
    fromSO => R1_inj_so,
    toCE => SIB_1_inj_toCE,
    toSE => SIB_1_inj_toSE,
    toUE => SIB_1_inj_toUE,
    toSEL => SIB_1_inj_toSEL,
    toRST => SIB_1_inj_toRST,
    toTCK => SIB_1_inj_toTCK,
    toSI => SIB_1_inj_toSI,
    fromF => '0',
    fromC => '1'
);
-- Router 1 checker status SIB
SIB_1_status : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_1_inj_so,
    CE => SIB_1_toCE,
    SE => SIB_1_toSE,
    UE => SIB_1_toUE,
    SEL => SIB_1_toSEL,
    RST => SIB_1_toRST,
    TCK => SIB_1_toTCK,
    SO => SIB_1_sta_so,
    toF => F_fromSIB_1_status,
    toC => C_fromSIB_1_status,
     -- Scan Interface  host ----------------
    fromSO => R1_sta_adapter_so,
    toCE => SIB_1_sta_toCE,
    toSE => SIB_1_sta_toSE,
    toUE => SIB_1_sta_toUE,
    toSEL => SIB_1_sta_toSEL,
    toRST => SIB_1_sta_toRST,
    toTCK => SIB_1_sta_toTCK,
    toSI => SIB_1_sta_toSI,
    fromF => F_R1,
    fromC => C_R1
);
-- Router 1 checker status IJTAG adapter
R1_status_adapter : AsyncDataRegisterAdapter
    generic map (Size => 25)
    port map (
    SI => SIB_1_sta_toSI,
    SO => R1_sta_adapter_so,
    SEL => SIB_1_sta_toSEL,
    ----------------------------------------     
    SE => SIB_1_sta_toSE,
    CE => SIB_1_sta_toCE,
    UE => SIB_1_sta_toUE,
    RST => SIB_1_sta_toRST,
    TCK => SIB_1_sta_toTCK,
      -- Data interface
    DI => R1_aggregated_fault_status,
    DO => R1_sta_adapter_do
);

R1_aggregated_fault_status <= link_faults_async_1 & turn_faults_async_1;
-----------------------------------
------ ROUTER 2 -------------------
-----------------------------------
-- Router R2 main SIB
SIB_2 : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_1_so,
    CE => SIB_main_toCE,
    SE => SIB_main_toSE,
    UE => SIB_main_toUE,
    SEL => SIB_main_toSEL,
    RST => SIB_main_toRST,
    TCK => SIB_main_toTCK,
    SO => SIB_2_so,
    toF => F_segtop_fromSIB_2,
    toC => C_segtop_fromSIB_2,
     -- Scan Interface  host ----------------
    fromSO => SIB_2_sta_so,
    toCE => SIB_2_toCE,
    toSE => SIB_2_toSE,
    toUE => SIB_2_toUE,
    toSEL => SIB_2_toSEL,
    toRST => SIB_2_toRST,
    toTCK => SIB_2_toTCK,
    toSI => SIB_2_toSI,
    fromF => toF_SIB_2,
    fromC => toC_SIB_2
);

toF_SIB_2 <= F_fromSIB_2_inj or  F_fromSIB_2_status;
toC_SIB_2 <= C_fromSIB_2_inj and C_fromSIB_2_status;

-- Router 2 fault injection SIB
SIB_2_injection : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_2_toSI,
    CE => SIB_2_toCE,
    SE => SIB_2_toSE,
    UE => SIB_2_toUE,
    SEL => SIB_2_toSEL,
    RST => SIB_2_toRST,
    TCK => SIB_2_toTCK,
    SO => SIB_2_inj_so,
    toF => F_fromSIB_2_inj,
    toC => C_fromSIB_2_inj,
     -- Scan Interface  host ----------------
    fromSO => R2_inj_so,
    toCE => SIB_2_inj_toCE,
    toSE => SIB_2_inj_toSE,
    toUE => SIB_2_inj_toUE,
    toSEL => SIB_2_inj_toSEL,
    toRST => SIB_2_inj_toRST,
    toTCK => SIB_2_inj_toTCK,
    toSI => SIB_2_inj_toSI,
    fromF => '0',
    fromC => '1'
);
-- Router 2 checker status SIB
SIB_2_status : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_2_inj_so,
    CE => SIB_2_toCE,
    SE => SIB_2_toSE,
    UE => SIB_2_toUE,
    SEL => SIB_2_toSEL,
    RST => SIB_2_toRST,
    TCK => SIB_2_toTCK,
    SO => SIB_2_sta_so,
    toF => F_fromSIB_2_status,
    toC => C_fromSIB_2_status,
     -- Scan Interface  host ----------------
    fromSO => R2_sta_adapter_so,
    toCE => SIB_2_sta_toCE,
    toSE => SIB_2_sta_toSE,
    toUE => SIB_2_sta_toUE,
    toSEL => SIB_2_sta_toSEL,
    toRST => SIB_2_sta_toRST,
    toTCK => SIB_2_sta_toTCK,
    toSI => SIB_2_sta_toSI,
    fromF => F_R2,
    fromC => C_R2
);
-- Router 2 checker status IJTAG adapter
R2_status_adapter : AsyncDataRegisterAdapter
    generic map (Size => 25)
    port map (
    SI => SIB_2_sta_toSI,
    SO => R2_sta_adapter_so,
    SEL => SIB_2_sta_toSEL,
    ----------------------------------------     
    SE => SIB_2_sta_toSE,
    CE => SIB_2_sta_toCE,
    UE => SIB_2_sta_toUE,
    RST => SIB_2_sta_toRST,
    TCK => SIB_2_sta_toTCK,
      -- Data interface
    DI => R2_aggregated_fault_status,
    DO => R2_sta_adapter_do
);

R2_aggregated_fault_status <= link_faults_async_2 & turn_faults_async_2;
-----------------------------------
------ ROUTER 3 -------------------
-----------------------------------
-- Router 3 main SIB
SIB_3 : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_2_so,
    CE => SIB_main_toCE,
    SE => SIB_main_toSE,
    UE => SIB_main_toUE,
    SEL => SIB_main_toSEL,
    RST => SIB_main_toRST,
    TCK => SIB_main_toTCK,
    SO => SIB_3_so,
    toF => F_segtop_fromSIB_3,
    toC => C_segtop_fromSIB_3,
     -- Scan Interface  host ----------------
    fromSO => SIB_3_sta_so,
    toCE => SIB_3_toCE,
    toSE => SIB_3_toSE,
    toUE => SIB_3_toUE,
    toSEL => SIB_3_toSEL,
    toRST => SIB_3_toRST,
    toTCK => SIB_3_toTCK,
    toSI => SIB_3_toSI,
    fromF => toF_SIB_3,
    fromC => toC_SIB_3
);

toF_SIB_3 <= F_fromSIB_3_inj or  F_fromSIB_3_status;
toC_SIB_3 <= C_fromSIB_3_inj and C_fromSIB_3_status;

-- Router 3 fault injection SIB
SIB_3_injection : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_3_toSI,
    CE => SIB_3_toCE,
    SE => SIB_3_toSE,
    UE => SIB_3_toUE,
    SEL => SIB_3_toSEL,
    RST => SIB_3_toRST,
    TCK => SIB_3_toTCK,
    SO => SIB_3_inj_so,
    toF => F_fromSIB_3_inj,
    toC => C_fromSIB_3_inj,
     -- Scan Interface  host ----------------
    fromSO => R3_inj_so,
    toCE => SIB_3_inj_toCE,
    toSE => SIB_3_inj_toSE,
    toUE => SIB_3_inj_toUE,
    toSEL => SIB_3_inj_toSEL,
    toRST => SIB_3_inj_toRST,
    toTCK => SIB_3_inj_toTCK,
    toSI => SIB_3_inj_toSI,
    fromF => '0',
    fromC => '1'
);
-- Router 3 checker status SIB
SIB_3_status : SIB_mux_pre_FCX_SELgate
    port map ( -- Scan Interface  client --------------
    SI => SIB_3_inj_so,
    CE => SIB_3_toCE,
    SE => SIB_3_toSE,
    UE => SIB_3_toUE,
    SEL => SIB_3_toSEL,
    RST => SIB_3_toRST,
    TCK => SIB_3_toTCK,
    SO => SIB_3_sta_so,
    toF => F_fromSIB_3_status,
    toC => C_fromSIB_3_status,
     -- Scan Interface  host ----------------
    fromSO => R3_sta_adapter_so,
    toCE => SIB_3_sta_toCE,
    toSE => SIB_3_sta_toSE,
    toUE => SIB_3_sta_toUE,
    toSEL => SIB_3_sta_toSEL,
    toRST => SIB_3_sta_toRST,
    toTCK => SIB_3_sta_toTCK,
    toSI => SIB_3_sta_toSI,
    fromF => F_R3,
    fromC => C_R3
);
-- Router 3 checker status IJTAG adapter
R3_status_adapter : AsyncDataRegisterAdapter
    generic map (Size => 25)
    port map (
    SI => SIB_3_sta_toSI,
    SO => R3_sta_adapter_so,
    SEL => SIB_3_sta_toSEL,
    ----------------------------------------     
    SE => SIB_3_sta_toSE,
    CE => SIB_3_sta_toCE,
    UE => SIB_3_sta_toUE,
    RST => SIB_3_sta_toRST,
    TCK => SIB_3_sta_toTCK,
      -- Data interface
    DI => R3_aggregated_fault_status,
    DO => R3_sta_adapter_do
);
    
R3_aggregated_fault_status <= link_faults_async_3 & turn_faults_async_3;

-- Fault flags are ORs of all fault signals coming from routers
F_R0 <= OR_REDUCE(link_faults_async_0&turn_faults_async_0);
F_R1 <= OR_REDUCE(link_faults_async_1&turn_faults_async_1);
F_R2 <= OR_REDUCE(link_faults_async_2&turn_faults_async_2);
F_R3 <= OR_REDUCE(link_faults_async_3&turn_faults_async_3);

-- A fault in a router does not need the whole system to be halted,
-- so lower priority fault can be used (F = 1, C = 1 in case of fault)
C_R0 <= '1';
C_R1 <= '1';
C_R2 <= '1';
C_R3 <= '1';

R_0: router_NW_credit_based_PD_C_SHMU 
    generic map (DATA_WIDTH =>DATA_WIDTH,         current_address => 0, Rxy_rst => 60,
        Cx_rst =>  10, NoC_size => 2, healthy_counter_threshold => 15, faulty_counter_threshold => 3, counter_depth => 4)
    port map(
    reset, clk,
	RX_E_0, RX_S_0, RX_L_0,
	credit_in_E_0, credit_in_S_0, credit_in_L_0,
	valid_in_E_0, valid_in_S_0, valid_in_L_0,
	valid_out_E_0, valid_out_S_0, valid_out_L_0,
	credit_out_E_0, credit_out_S_0, credit_out_L_0,
	TX_E_0, TX_S_0, TX_L_0,
	Faulty_E_in0,Faulty_S_in0,
	Faulty_E_out0,Faulty_S_out0,
	-- should be connected to NI
	link_faults_0, turn_faults_0,
	Rxy_reconf_PE_0, Cx_reconf_PE_0, Reconfig_command_0, 
	-- fault injector shift register with serial input signals
    SIB_0_inj_toTCK, SIB_0_inj_toSE, SIB_0_inj_toUE, SIB_0_inj_toSI, R0_inj_so,
    -- the non-classified fault information
    link_faults_async_0, turn_faults_async_0
 ); 

R_1: router_NE_credit_based_PD_C_SHMU 
    generic map (DATA_WIDTH =>DATA_WIDTH,         current_address => 1, Rxy_rst => 60,
        Cx_rst =>  12, NoC_size => 2, healthy_counter_threshold => 15, faulty_counter_threshold => 3, counter_depth => 4)
    port map(
    reset, clk,
	RX_W_1, RX_S_1, RX_L_1,
	credit_in_W_1, credit_in_S_1, credit_in_L_1,
	valid_in_W_1, valid_in_S_1, valid_in_L_1,
	valid_out_W_1, valid_out_S_1, valid_out_L_1,
	credit_out_W_1, credit_out_S_1, credit_out_L_1,
	TX_W_1, TX_S_1, TX_L_1,
	Faulty_W_in1,Faulty_S_in1,
	Faulty_W_out1,Faulty_S_out1,
	-- should be connected to NI
	link_faults_1, turn_faults_1,
	Rxy_reconf_PE_1, Cx_reconf_PE_1, Reconfig_command_1, 
    -- fault injector shift register with serial input signals
    SIB_1_inj_toTCK, SIB_1_inj_toSE, SIB_1_inj_toUE, SIB_1_inj_toSI, R1_inj_so,
    -- the non-classified fault information
    link_faults_async_1, turn_faults_async_1
 ); 
    
R_2: router_SW_credit_based_PD_C_SHMU 
    generic map (DATA_WIDTH =>DATA_WIDTH,         current_address => 2, Rxy_rst => 60,
        Cx_rst =>  3, NoC_size => 2, healthy_counter_threshold => 15, faulty_counter_threshold => 3, counter_depth => 4)
    port map(
    reset, clk,
	RX_N_2, RX_E_2, RX_L_2,
	credit_in_N_2, credit_in_E_2, credit_in_L_2,
	valid_in_N_2, valid_in_E_2, valid_in_L_2,
	valid_out_N_2, valid_out_E_2, valid_out_L_2,
	credit_out_N_2, credit_out_E_2, credit_out_L_2,
	TX_N_2, TX_E_2, TX_L_2,
	Faulty_N_in2,Faulty_E_in2,
	Faulty_N_out2,Faulty_E_out2,
	-- should be connected to NI
	link_faults_2, turn_faults_2,
	Rxy_reconf_PE_2, Cx_reconf_PE_2, Reconfig_command_2, 
    -- fault injector shift register with serial input signals
    SIB_2_inj_toTCK, SIB_2_inj_toSE, SIB_2_inj_toUE, SIB_2_inj_toSI, R2_inj_so,
    -- the non-classified fault information
    link_faults_async_2, turn_faults_async_2
 ); 

R_3: router_SE_credit_based_PD_C_SHMU 
    generic map (DATA_WIDTH =>DATA_WIDTH,         current_address => 3, Rxy_rst => 60,
        Cx_rst =>  5, NoC_size => 2, healthy_counter_threshold => 15, faulty_counter_threshold => 3, counter_depth => 4)
    port map(
    reset, clk,
	RX_N_3, RX_W_3, RX_L_3,
	credit_in_N_3, credit_in_W_3, credit_in_L_3,
	valid_in_N_3, valid_in_W_3, valid_in_L_3,
	valid_out_N_3, valid_out_W_3, valid_out_L_3,
	credit_out_N_3, credit_out_W_3, credit_out_L_3,
	TX_N_3, TX_W_3, TX_L_3,
	Faulty_N_in3,Faulty_W_in3,
	Faulty_N_out3,Faulty_W_out3,
	-- should be connected to NI
	link_faults_3, turn_faults_3,
	Rxy_reconf_PE_3, Cx_reconf_PE_3, Reconfig_command_3, 
    -- fault injector shift register with serial input signals
    SIB_3_inj_toTCK, SIB_3_inj_toSE, SIB_3_inj_toUE, SIB_3_inj_toSI, R3_inj_so, 
    -- the non-classified fault information
    link_faults_async_3, turn_faults_async_3
 ); 

---------------------------------------------------------------
-- binding the routers together
-- vertical ins/outs
-- connecting router: 0 to router: 2 and vice versa
RX_N_2<= TX_S_0;
RX_S_0<= TX_N_2;
-------------------
-- connecting router: 1 to router: 3 and vice versa
RX_N_3<= TX_S_1;
RX_S_1<= TX_N_3;
-------------------

-- horizontal ins/outs
-- connecting router: 0 to router: 1 and vice versa
RX_E_0 <= TX_W_1;
RX_W_1 <= TX_E_0;
-------------------
-- connecting router: 2 to router: 3 and vice versa
RX_E_2 <= TX_W_3;
RX_W_3 <= TX_E_2;
-------------------
---------------------------------------------------------------
-- binding the routers together
-- connecting router: 0 to router: 2 and vice versa
valid_in_N_2 <= valid_out_S_0;
valid_in_S_0 <= valid_out_N_2;
credit_in_S_0 <= credit_out_N_2;
credit_in_N_2 <= credit_out_S_0;
-------------------
-- connecting router: 1 to router: 3 and vice versa
valid_in_N_3 <= valid_out_S_1;
valid_in_S_1 <= valid_out_N_3;
credit_in_S_1 <= credit_out_N_3;
credit_in_N_3 <= credit_out_S_1;
-------------------

-- connecting router: 0 to router: 1 and vice versa
valid_in_E_0 <= valid_out_W_1;
valid_in_W_1 <= valid_out_E_0;
credit_in_W_1 <= credit_out_E_0;
credit_in_E_0 <= credit_out_W_1;
-------------------
-- connecting router: 2 to router: 3 and vice versa
valid_in_E_2 <= valid_out_W_3;
valid_in_W_3 <= valid_out_E_2;
credit_in_W_3 <= credit_out_E_2;
credit_in_E_2 <= credit_out_W_3;
-------------------
Faulty_S_in0 <= Faulty_N_out2;
Faulty_E_in0 <= Faulty_W_out1;
Faulty_S_in1 <= Faulty_N_out3;
Faulty_W_in1 <= Faulty_E_out0;
Faulty_N_in2 <= Faulty_S_out0;
Faulty_E_in2 <= Faulty_W_out3;
Faulty_N_in3 <= Faulty_S_out1;
Faulty_W_in3 <= Faulty_E_out2;
end;
